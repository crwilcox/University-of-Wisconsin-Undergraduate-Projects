
module Packet_Queue_0 ( Clk_r, Rst_n, Packet_In, Read_Ack, Write_Ack, 
        Packet_Out, Empty, Full );
  input [31:0] Packet_In;
  output [31:0] Packet_Out;
  input Clk_r, Rst_n, Read_Ack, Write_Ack;
  output Empty, Full;
  wire   \Queue[4][31] , \Queue[4][30] , \Queue[4][29] , \Queue[4][28] ,
         \Queue[4][27] , \Queue[4][26] , \Queue[4][25] , \Queue[4][24] ,
         \Queue[4][23] , \Queue[4][22] , \Queue[4][21] , \Queue[4][20] ,
         \Queue[4][19] , \Queue[4][18] , \Queue[4][17] , \Queue[4][16] ,
         \Queue[4][15] , \Queue[4][14] , \Queue[4][13] , \Queue[4][12] ,
         \Queue[4][11] , \Queue[4][10] , \Queue[4][9] , \Queue[4][8] ,
         \Queue[4][7] , \Queue[4][6] , \Queue[4][5] , \Queue[4][4] ,
         \Queue[4][3] , \Queue[4][2] , \Queue[4][1] , \Queue[4][0] ,
         \Queue[3][31] , \Queue[3][30] , \Queue[3][29] , \Queue[3][28] ,
         \Queue[3][27] , \Queue[3][26] , \Queue[3][25] , \Queue[3][24] ,
         \Queue[3][23] , \Queue[3][22] , \Queue[3][21] , \Queue[3][20] ,
         \Queue[3][19] , \Queue[3][18] , \Queue[3][17] , \Queue[3][16] ,
         \Queue[3][15] , \Queue[3][14] , \Queue[3][13] , \Queue[3][12] ,
         \Queue[3][11] , \Queue[3][10] , \Queue[3][9] , \Queue[3][8] ,
         \Queue[3][7] , \Queue[3][6] , \Queue[3][5] , \Queue[3][4] ,
         \Queue[3][3] , \Queue[3][2] , \Queue[3][1] , \Queue[3][0] ,
         \Queue[2][31] , \Queue[2][30] , \Queue[2][29] , \Queue[2][28] ,
         \Queue[2][27] , \Queue[2][26] , \Queue[2][25] , \Queue[2][24] ,
         \Queue[2][23] , \Queue[2][22] , \Queue[2][21] , \Queue[2][20] ,
         \Queue[2][19] , \Queue[2][18] , \Queue[2][17] , \Queue[2][16] ,
         \Queue[2][15] , \Queue[2][14] , \Queue[2][13] , \Queue[2][12] ,
         \Queue[2][11] , \Queue[2][10] , \Queue[2][9] , \Queue[2][8] ,
         \Queue[2][7] , \Queue[2][6] , \Queue[2][5] , \Queue[2][4] ,
         \Queue[2][3] , \Queue[2][2] , \Queue[2][1] , \Queue[2][0] ,
         \Queue[1][31] , \Queue[1][30] , \Queue[1][29] , \Queue[1][28] ,
         \Queue[1][27] , \Queue[1][26] , \Queue[1][25] , \Queue[1][24] ,
         \Queue[1][23] , \Queue[1][22] , \Queue[1][21] , \Queue[1][20] ,
         \Queue[1][19] , \Queue[1][18] , \Queue[1][17] , \Queue[1][16] ,
         \Queue[1][15] , \Queue[1][14] , \Queue[1][13] , \Queue[1][12] ,
         \Queue[1][11] , \Queue[1][10] , \Queue[1][9] , \Queue[1][8] ,
         \Queue[1][7] , \Queue[1][6] , \Queue[1][5] , \Queue[1][4] ,
         \Queue[1][3] , \Queue[1][2] , \Queue[1][1] , \Queue[1][0] , n1, n2,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n373, n374, n375, n376,
         n377, n378, n379;
  wire   [2:0] Count;

  FDN2QM1P \Count_reg[0]  ( .D(n372), .CPN(Clk_r), .CD(Rst_n), .Q(Count[0]) );
  FDN2QM1P \Count_reg[1]  ( .D(n371), .CPN(Clk_r), .CD(Rst_n), .Q(Count[1]) );
  FDN2QM1P \Count_reg[2]  ( .D(n370), .CPN(Clk_r), .CD(Rst_n), .Q(Count[2]) );
  FDN1QM1P \Queue_reg[4][30]  ( .D(n338), .CPN(Clk_r), .Q(\Queue[4][30] ) );
  FDN1QM1P \Queue_reg[3][30]  ( .D(n210), .CPN(Clk_r), .Q(\Queue[3][30] ) );
  FDN1QM1P \Queue_reg[2][30]  ( .D(n242), .CPN(Clk_r), .Q(\Queue[2][30] ) );
  FDN1QM1P \Queue_reg[4][29]  ( .D(n339), .CPN(Clk_r), .Q(\Queue[4][29] ) );
  FDN1QM1P \Queue_reg[3][29]  ( .D(n211), .CPN(Clk_r), .Q(\Queue[3][29] ) );
  FDN1QM1P \Queue_reg[2][29]  ( .D(n243), .CPN(Clk_r), .Q(\Queue[2][29] ) );
  FDN1QM1P \Queue_reg[4][28]  ( .D(n340), .CPN(Clk_r), .Q(\Queue[4][28] ) );
  FDN1QM1P \Queue_reg[3][28]  ( .D(n212), .CPN(Clk_r), .Q(\Queue[3][28] ) );
  FDN1QM1P \Queue_reg[2][28]  ( .D(n244), .CPN(Clk_r), .Q(\Queue[2][28] ) );
  FDN1QM1P \Queue_reg[4][27]  ( .D(n341), .CPN(Clk_r), .Q(\Queue[4][27] ) );
  FDN1QM1P \Queue_reg[3][27]  ( .D(n213), .CPN(Clk_r), .Q(\Queue[3][27] ) );
  FDN1QM1P \Queue_reg[2][27]  ( .D(n245), .CPN(Clk_r), .Q(\Queue[2][27] ) );
  FDN1QM1P \Queue_reg[4][26]  ( .D(n342), .CPN(Clk_r), .Q(\Queue[4][26] ) );
  FDN1QM1P \Queue_reg[3][26]  ( .D(n214), .CPN(Clk_r), .Q(\Queue[3][26] ) );
  FDN1QM1P \Queue_reg[2][26]  ( .D(n246), .CPN(Clk_r), .Q(\Queue[2][26] ) );
  FDN1QM1P \Queue_reg[4][25]  ( .D(n343), .CPN(Clk_r), .Q(\Queue[4][25] ) );
  FDN1QM1P \Queue_reg[3][25]  ( .D(n215), .CPN(Clk_r), .Q(\Queue[3][25] ) );
  FDN1QM1P \Queue_reg[2][25]  ( .D(n247), .CPN(Clk_r), .Q(\Queue[2][25] ) );
  FDN1QM1P \Queue_reg[4][24]  ( .D(n344), .CPN(Clk_r), .Q(\Queue[4][24] ) );
  FDN1QM1P \Queue_reg[3][24]  ( .D(n216), .CPN(Clk_r), .Q(\Queue[3][24] ) );
  FDN1QM1P \Queue_reg[2][24]  ( .D(n248), .CPN(Clk_r), .Q(\Queue[2][24] ) );
  FDN1QM1P \Queue_reg[4][23]  ( .D(n345), .CPN(Clk_r), .Q(\Queue[4][23] ) );
  FDN1QM1P \Queue_reg[3][23]  ( .D(n217), .CPN(Clk_r), .Q(\Queue[3][23] ) );
  FDN1QM1P \Queue_reg[2][23]  ( .D(n249), .CPN(Clk_r), .Q(\Queue[2][23] ) );
  FDN1QM1P \Queue_reg[4][22]  ( .D(n346), .CPN(Clk_r), .Q(\Queue[4][22] ) );
  FDN1QM1P \Queue_reg[3][22]  ( .D(n218), .CPN(Clk_r), .Q(\Queue[3][22] ) );
  FDN1QM1P \Queue_reg[2][22]  ( .D(n250), .CPN(Clk_r), .Q(\Queue[2][22] ) );
  FDN1QM1P \Queue_reg[4][21]  ( .D(n347), .CPN(Clk_r), .Q(\Queue[4][21] ) );
  FDN1QM1P \Queue_reg[3][21]  ( .D(n219), .CPN(Clk_r), .Q(\Queue[3][21] ) );
  FDN1QM1P \Queue_reg[2][21]  ( .D(n251), .CPN(Clk_r), .Q(\Queue[2][21] ) );
  FDN1QM1P \Queue_reg[4][20]  ( .D(n348), .CPN(Clk_r), .Q(\Queue[4][20] ) );
  FDN1QM1P \Queue_reg[3][20]  ( .D(n220), .CPN(Clk_r), .Q(\Queue[3][20] ) );
  FDN1QM1P \Queue_reg[2][20]  ( .D(n252), .CPN(Clk_r), .Q(\Queue[2][20] ) );
  FDN1QM1P \Queue_reg[4][19]  ( .D(n349), .CPN(Clk_r), .Q(\Queue[4][19] ) );
  FDN1QM1P \Queue_reg[3][19]  ( .D(n221), .CPN(Clk_r), .Q(\Queue[3][19] ) );
  FDN1QM1P \Queue_reg[2][19]  ( .D(n253), .CPN(Clk_r), .Q(\Queue[2][19] ) );
  FDN1QM1P \Queue_reg[4][18]  ( .D(n350), .CPN(Clk_r), .Q(\Queue[4][18] ) );
  FDN1QM1P \Queue_reg[3][18]  ( .D(n222), .CPN(Clk_r), .Q(\Queue[3][18] ) );
  FDN1QM1P \Queue_reg[2][18]  ( .D(n254), .CPN(Clk_r), .Q(\Queue[2][18] ) );
  FDN1QM1P \Queue_reg[4][17]  ( .D(n351), .CPN(Clk_r), .Q(\Queue[4][17] ) );
  FDN1QM1P \Queue_reg[3][17]  ( .D(n223), .CPN(Clk_r), .Q(\Queue[3][17] ) );
  FDN1QM1P \Queue_reg[2][17]  ( .D(n255), .CPN(Clk_r), .Q(\Queue[2][17] ) );
  FDN1QM1P \Queue_reg[4][16]  ( .D(n352), .CPN(Clk_r), .Q(\Queue[4][16] ) );
  FDN1QM1P \Queue_reg[3][16]  ( .D(n224), .CPN(Clk_r), .Q(\Queue[3][16] ) );
  FDN1QM1P \Queue_reg[2][16]  ( .D(n256), .CPN(Clk_r), .Q(\Queue[2][16] ) );
  FDN1QM1P \Queue_reg[4][15]  ( .D(n353), .CPN(Clk_r), .Q(\Queue[4][15] ) );
  FDN1QM1P \Queue_reg[3][15]  ( .D(n225), .CPN(Clk_r), .Q(\Queue[3][15] ) );
  FDN1QM1P \Queue_reg[2][15]  ( .D(n257), .CPN(Clk_r), .Q(\Queue[2][15] ) );
  FDN1QM1P \Queue_reg[4][14]  ( .D(n354), .CPN(Clk_r), .Q(\Queue[4][14] ) );
  FDN1QM1P \Queue_reg[3][14]  ( .D(n226), .CPN(Clk_r), .Q(\Queue[3][14] ) );
  FDN1QM1P \Queue_reg[2][14]  ( .D(n258), .CPN(Clk_r), .Q(\Queue[2][14] ) );
  FDN1QM1P \Queue_reg[4][13]  ( .D(n355), .CPN(Clk_r), .Q(\Queue[4][13] ) );
  FDN1QM1P \Queue_reg[3][13]  ( .D(n227), .CPN(Clk_r), .Q(\Queue[3][13] ) );
  FDN1QM1P \Queue_reg[2][13]  ( .D(n259), .CPN(Clk_r), .Q(\Queue[2][13] ) );
  FDN1QM1P \Queue_reg[4][12]  ( .D(n356), .CPN(Clk_r), .Q(\Queue[4][12] ) );
  FDN1QM1P \Queue_reg[3][12]  ( .D(n228), .CPN(Clk_r), .Q(\Queue[3][12] ) );
  FDN1QM1P \Queue_reg[2][12]  ( .D(n260), .CPN(Clk_r), .Q(\Queue[2][12] ) );
  FDN1QM1P \Queue_reg[4][11]  ( .D(n357), .CPN(Clk_r), .Q(\Queue[4][11] ) );
  FDN1QM1P \Queue_reg[3][11]  ( .D(n229), .CPN(Clk_r), .Q(\Queue[3][11] ) );
  FDN1QM1P \Queue_reg[2][11]  ( .D(n261), .CPN(Clk_r), .Q(\Queue[2][11] ) );
  FDN1QM1P \Queue_reg[4][10]  ( .D(n358), .CPN(Clk_r), .Q(\Queue[4][10] ) );
  FDN1QM1P \Queue_reg[3][10]  ( .D(n230), .CPN(Clk_r), .Q(\Queue[3][10] ) );
  FDN1QM1P \Queue_reg[2][10]  ( .D(n262), .CPN(Clk_r), .Q(\Queue[2][10] ) );
  FDN1QM1P \Queue_reg[4][9]  ( .D(n359), .CPN(Clk_r), .Q(\Queue[4][9] ) );
  FDN1QM1P \Queue_reg[3][9]  ( .D(n231), .CPN(Clk_r), .Q(\Queue[3][9] ) );
  FDN1QM1P \Queue_reg[2][9]  ( .D(n263), .CPN(Clk_r), .Q(\Queue[2][9] ) );
  FDN1QM1P \Queue_reg[4][8]  ( .D(n360), .CPN(Clk_r), .Q(\Queue[4][8] ) );
  FDN1QM1P \Queue_reg[3][8]  ( .D(n232), .CPN(Clk_r), .Q(\Queue[3][8] ) );
  FDN1QM1P \Queue_reg[2][8]  ( .D(n264), .CPN(Clk_r), .Q(\Queue[2][8] ) );
  FDN1QM1P \Queue_reg[4][7]  ( .D(n361), .CPN(Clk_r), .Q(\Queue[4][7] ) );
  FDN1QM1P \Queue_reg[3][7]  ( .D(n233), .CPN(Clk_r), .Q(\Queue[3][7] ) );
  FDN1QM1P \Queue_reg[2][7]  ( .D(n265), .CPN(Clk_r), .Q(\Queue[2][7] ) );
  FDN1QM1P \Queue_reg[4][6]  ( .D(n362), .CPN(Clk_r), .Q(\Queue[4][6] ) );
  FDN1QM1P \Queue_reg[3][6]  ( .D(n234), .CPN(Clk_r), .Q(\Queue[3][6] ) );
  FDN1QM1P \Queue_reg[2][6]  ( .D(n266), .CPN(Clk_r), .Q(\Queue[2][6] ) );
  FDN1QM1P \Queue_reg[4][5]  ( .D(n363), .CPN(Clk_r), .Q(\Queue[4][5] ) );
  FDN1QM1P \Queue_reg[3][5]  ( .D(n235), .CPN(Clk_r), .Q(\Queue[3][5] ) );
  FDN1QM1P \Queue_reg[2][5]  ( .D(n267), .CPN(Clk_r), .Q(\Queue[2][5] ) );
  FDN1QM1P \Queue_reg[4][4]  ( .D(n364), .CPN(Clk_r), .Q(\Queue[4][4] ) );
  FDN1QM1P \Queue_reg[3][4]  ( .D(n236), .CPN(Clk_r), .Q(\Queue[3][4] ) );
  FDN1QM1P \Queue_reg[2][4]  ( .D(n268), .CPN(Clk_r), .Q(\Queue[2][4] ) );
  FDN1QM1P \Queue_reg[4][3]  ( .D(n365), .CPN(Clk_r), .Q(\Queue[4][3] ) );
  FDN1QM1P \Queue_reg[3][3]  ( .D(n237), .CPN(Clk_r), .Q(\Queue[3][3] ) );
  FDN1QM1P \Queue_reg[2][3]  ( .D(n269), .CPN(Clk_r), .Q(\Queue[2][3] ) );
  FDN1QM1P \Queue_reg[4][2]  ( .D(n366), .CPN(Clk_r), .Q(\Queue[4][2] ) );
  FDN1QM1P \Queue_reg[3][2]  ( .D(n238), .CPN(Clk_r), .Q(\Queue[3][2] ) );
  FDN1QM1P \Queue_reg[2][2]  ( .D(n270), .CPN(Clk_r), .Q(\Queue[2][2] ) );
  FDN1QM1P \Queue_reg[4][1]  ( .D(n367), .CPN(Clk_r), .Q(\Queue[4][1] ) );
  FDN1QM1P \Queue_reg[3][1]  ( .D(n239), .CPN(Clk_r), .Q(\Queue[3][1] ) );
  FDN1QM1P \Queue_reg[2][1]  ( .D(n271), .CPN(Clk_r), .Q(\Queue[2][1] ) );
  FDN1QM1P \Queue_reg[4][0]  ( .D(n368), .CPN(Clk_r), .Q(\Queue[4][0] ) );
  FDN1QM1P \Queue_reg[3][0]  ( .D(n240), .CPN(Clk_r), .Q(\Queue[3][0] ) );
  FDN1QM1P \Queue_reg[2][0]  ( .D(n272), .CPN(Clk_r), .Q(\Queue[2][0] ) );
  FDN1QM1P \Queue_reg[4][31]  ( .D(n369), .CPN(Clk_r), .Q(\Queue[4][31] ) );
  FDN1QM1P \Queue_reg[3][31]  ( .D(n209), .CPN(Clk_r), .Q(\Queue[3][31] ) );
  FDN1QM1P \Queue_reg[2][31]  ( .D(n241), .CPN(Clk_r), .Q(\Queue[2][31] ) );
  FDN2QM1P Full_reg ( .D(n337), .CPN(Clk_r), .CD(Rst_n), .Q(Full) );
  FDN1QM1P \Queue_reg[1][31]  ( .D(n305), .CPN(Clk_r), .Q(\Queue[1][31] ) );
  FDN1QM1P \Queue_reg[0][31]  ( .D(n273), .CPN(Clk_r), .Q(Packet_Out[31]) );
  FDN1QM1P \Queue_reg[1][30]  ( .D(n306), .CPN(Clk_r), .Q(\Queue[1][30] ) );
  FDN1QM1P \Queue_reg[0][30]  ( .D(n274), .CPN(Clk_r), .Q(Packet_Out[30]) );
  FDN1QM1P \Queue_reg[1][29]  ( .D(n307), .CPN(Clk_r), .Q(\Queue[1][29] ) );
  FDN1QM1P \Queue_reg[0][29]  ( .D(n275), .CPN(Clk_r), .Q(Packet_Out[29]) );
  FDN1QM1P \Queue_reg[1][28]  ( .D(n308), .CPN(Clk_r), .Q(\Queue[1][28] ) );
  FDN1QM1P \Queue_reg[0][28]  ( .D(n276), .CPN(Clk_r), .Q(Packet_Out[28]) );
  FDN1QM1P \Queue_reg[1][27]  ( .D(n309), .CPN(Clk_r), .Q(\Queue[1][27] ) );
  FDN1QM1P \Queue_reg[0][27]  ( .D(n277), .CPN(Clk_r), .Q(Packet_Out[27]) );
  FDN1QM1P \Queue_reg[1][26]  ( .D(n310), .CPN(Clk_r), .Q(\Queue[1][26] ) );
  FDN1QM1P \Queue_reg[0][26]  ( .D(n278), .CPN(Clk_r), .Q(Packet_Out[26]) );
  FDN1QM1P \Queue_reg[1][25]  ( .D(n311), .CPN(Clk_r), .Q(\Queue[1][25] ) );
  FDN1QM1P \Queue_reg[0][25]  ( .D(n279), .CPN(Clk_r), .Q(Packet_Out[25]) );
  FDN1QM1P \Queue_reg[1][24]  ( .D(n312), .CPN(Clk_r), .Q(\Queue[1][24] ) );
  FDN1QM1P \Queue_reg[0][24]  ( .D(n280), .CPN(Clk_r), .Q(Packet_Out[24]) );
  FDN1QM1P \Queue_reg[1][23]  ( .D(n313), .CPN(Clk_r), .Q(\Queue[1][23] ) );
  FDN1QM1P \Queue_reg[0][23]  ( .D(n281), .CPN(Clk_r), .Q(Packet_Out[23]) );
  FDN1QM1P \Queue_reg[1][22]  ( .D(n314), .CPN(Clk_r), .Q(\Queue[1][22] ) );
  FDN1QM1P \Queue_reg[0][22]  ( .D(n282), .CPN(Clk_r), .Q(Packet_Out[22]) );
  FDN1QM1P \Queue_reg[1][21]  ( .D(n315), .CPN(Clk_r), .Q(\Queue[1][21] ) );
  FDN1QM1P \Queue_reg[0][21]  ( .D(n283), .CPN(Clk_r), .Q(Packet_Out[21]) );
  FDN1QM1P \Queue_reg[1][20]  ( .D(n316), .CPN(Clk_r), .Q(\Queue[1][20] ) );
  FDN1QM1P \Queue_reg[0][20]  ( .D(n284), .CPN(Clk_r), .Q(Packet_Out[20]) );
  FDN1QM1P \Queue_reg[1][19]  ( .D(n317), .CPN(Clk_r), .Q(\Queue[1][19] ) );
  FDN1QM1P \Queue_reg[0][19]  ( .D(n285), .CPN(Clk_r), .Q(Packet_Out[19]) );
  FDN1QM1P \Queue_reg[1][18]  ( .D(n318), .CPN(Clk_r), .Q(\Queue[1][18] ) );
  FDN1QM1P \Queue_reg[0][18]  ( .D(n286), .CPN(Clk_r), .Q(Packet_Out[18]) );
  FDN1QM1P \Queue_reg[1][17]  ( .D(n319), .CPN(Clk_r), .Q(\Queue[1][17] ) );
  FDN1QM1P \Queue_reg[0][17]  ( .D(n287), .CPN(Clk_r), .Q(Packet_Out[17]) );
  FDN1QM1P \Queue_reg[1][16]  ( .D(n320), .CPN(Clk_r), .Q(\Queue[1][16] ) );
  FDN1QM1P \Queue_reg[0][16]  ( .D(n288), .CPN(Clk_r), .Q(Packet_Out[16]) );
  FDN1QM1P \Queue_reg[1][15]  ( .D(n321), .CPN(Clk_r), .Q(\Queue[1][15] ) );
  FDN1QM1P \Queue_reg[0][15]  ( .D(n289), .CPN(Clk_r), .Q(Packet_Out[15]) );
  FDN1QM1P \Queue_reg[1][14]  ( .D(n322), .CPN(Clk_r), .Q(\Queue[1][14] ) );
  FDN1QM1P \Queue_reg[0][14]  ( .D(n290), .CPN(Clk_r), .Q(Packet_Out[14]) );
  FDN1QM1P \Queue_reg[1][13]  ( .D(n323), .CPN(Clk_r), .Q(\Queue[1][13] ) );
  FDN1QM1P \Queue_reg[0][13]  ( .D(n291), .CPN(Clk_r), .Q(Packet_Out[13]) );
  FDN1QM1P \Queue_reg[1][12]  ( .D(n324), .CPN(Clk_r), .Q(\Queue[1][12] ) );
  FDN1QM1P \Queue_reg[0][12]  ( .D(n292), .CPN(Clk_r), .Q(Packet_Out[12]) );
  FDN1QM1P \Queue_reg[1][11]  ( .D(n325), .CPN(Clk_r), .Q(\Queue[1][11] ) );
  FDN1QM1P \Queue_reg[0][11]  ( .D(n293), .CPN(Clk_r), .Q(Packet_Out[11]) );
  FDN1QM1P \Queue_reg[1][10]  ( .D(n326), .CPN(Clk_r), .Q(\Queue[1][10] ) );
  FDN1QM1P \Queue_reg[0][10]  ( .D(n294), .CPN(Clk_r), .Q(Packet_Out[10]) );
  FDN1QM1P \Queue_reg[1][9]  ( .D(n327), .CPN(Clk_r), .Q(\Queue[1][9] ) );
  FDN1QM1P \Queue_reg[0][9]  ( .D(n295), .CPN(Clk_r), .Q(Packet_Out[9]) );
  FDN1QM1P \Queue_reg[1][8]  ( .D(n328), .CPN(Clk_r), .Q(\Queue[1][8] ) );
  FDN1QM1P \Queue_reg[0][8]  ( .D(n296), .CPN(Clk_r), .Q(Packet_Out[8]) );
  FDN1QM1P \Queue_reg[1][7]  ( .D(n329), .CPN(Clk_r), .Q(\Queue[1][7] ) );
  FDN1QM1P \Queue_reg[0][7]  ( .D(n297), .CPN(Clk_r), .Q(Packet_Out[7]) );
  FDN1QM1P \Queue_reg[1][6]  ( .D(n330), .CPN(Clk_r), .Q(\Queue[1][6] ) );
  FDN1QM1P \Queue_reg[0][6]  ( .D(n298), .CPN(Clk_r), .Q(Packet_Out[6]) );
  FDN1QM1P \Queue_reg[1][5]  ( .D(n331), .CPN(Clk_r), .Q(\Queue[1][5] ) );
  FDN1QM1P \Queue_reg[0][5]  ( .D(n299), .CPN(Clk_r), .Q(Packet_Out[5]) );
  FDN1QM1P \Queue_reg[1][4]  ( .D(n332), .CPN(Clk_r), .Q(\Queue[1][4] ) );
  FDN1QM1P \Queue_reg[0][4]  ( .D(n300), .CPN(Clk_r), .Q(Packet_Out[4]) );
  FDN1QM1P \Queue_reg[1][3]  ( .D(n333), .CPN(Clk_r), .Q(\Queue[1][3] ) );
  FDN1QM1P \Queue_reg[0][3]  ( .D(n301), .CPN(Clk_r), .Q(Packet_Out[3]) );
  FDN1QM1P \Queue_reg[1][2]  ( .D(n334), .CPN(Clk_r), .Q(\Queue[1][2] ) );
  FDN1QM1P \Queue_reg[0][2]  ( .D(n302), .CPN(Clk_r), .Q(Packet_Out[2]) );
  FDN1QM1P \Queue_reg[1][1]  ( .D(n335), .CPN(Clk_r), .Q(\Queue[1][1] ) );
  FDN1QM1P \Queue_reg[0][1]  ( .D(n303), .CPN(Clk_r), .Q(Packet_Out[1]) );
  FDN1QM1P \Queue_reg[1][0]  ( .D(n336), .CPN(Clk_r), .Q(\Queue[1][0] ) );
  FDN1QM1P \Queue_reg[0][0]  ( .D(n304), .CPN(Clk_r), .Q(Packet_Out[0]) );
  FDN2QM1P Empty_reg ( .D(n1), .CPN(Clk_r), .CD(Rst_n), .Q(n2) );
  ND2M1P U3 ( .A(Read_Ack), .B(Rst_n), .Z(n144) );
  N1M1P U4 ( .A(Read_Ack), .Z(n140) );
  N1M1P U5 ( .A(n3), .Z(n102) );
  OAI211M4P U6 ( .A(n103), .B(n140), .C(n3), .D(n27), .Z(n62) );
  AOI21M3P U7 ( .A(n3), .B(n143), .C(n144), .Z(n135) );
  OAI211M4P U8 ( .A(n143), .B(n140), .C(n3), .D(n101), .Z(n138) );
  OAI211M4P U9 ( .A(n145), .B(n140), .C(n3), .D(n139), .Z(n375) );
  NR2I1M8P U10 ( .A(n64), .B(n24), .Z(n23) );
  AOI21M3P U11 ( .A(n3), .B(n103), .C(n144), .Z(n60) );
  AOI21M3P U12 ( .A(n3), .B(n145), .C(n144), .Z(n208) );
  AOI21M3P U13 ( .A(n3), .B(n379), .C(n144), .Z(n98) );
  NR3M1P U14 ( .A(Count[2]), .B(n26), .C(n25), .Z(n143) );
  BUFM6P U15 ( .A(Write_Ack), .Z(n3) );
  BUFM3P U16 ( .A(n100), .Z(n10) );
  OAI211M2P U17 ( .A(n103), .B(n142), .C(Rst_n), .D(n141), .Z(n136) );
  OAI211M2P U18 ( .A(n143), .B(n142), .C(Rst_n), .D(n141), .Z(n373) );
  ND2M1P U19 ( .A(n21), .B(Rst_n), .Z(n64) );
  N1M1P U20 ( .A(n145), .Z(n24) );
  NR2M2P U21 ( .A(Read_Ack), .B(n102), .Z(n21) );
  NR3M1P U22 ( .A(Count[0]), .B(Count[1]), .C(n22), .Z(n145) );
  NR3M1P U23 ( .A(Count[0]), .B(Count[2]), .C(n25), .Z(n103) );
  NR3M1P U24 ( .A(n26), .B(Count[2]), .C(Count[1]), .Z(n379) );
  N1M1P U25 ( .A(Count[2]), .Z(n22) );
  N1M1P U26 ( .A(Count[1]), .Z(n25) );
  N1M1P U27 ( .A(Count[0]), .Z(n26) );
  N1M1P U28 ( .A(Packet_In[25]), .Z(n197) );
  N1M1P U29 ( .A(Packet_In[26]), .Z(n199) );
  N1M1P U30 ( .A(Packet_In[23]), .Z(n193) );
  N1M1P U31 ( .A(Packet_In[29]), .Z(n205) );
  N1M1P U32 ( .A(Packet_In[31]), .Z(n376) );
  N1M1P U33 ( .A(Packet_In[28]), .Z(n203) );
  N1M1P U34 ( .A(Packet_In[27]), .Z(n201) );
  N1M1P U35 ( .A(Packet_In[24]), .Z(n195) );
  N1M1P U36 ( .A(Packet_In[22]), .Z(n191) );
  N1M1P U37 ( .A(Packet_In[20]), .Z(n187) );
  N1M1P U38 ( .A(Packet_In[21]), .Z(n189) );
  N1M1P U39 ( .A(Packet_In[12]), .Z(n171) );
  N1M1P U40 ( .A(Packet_In[10]), .Z(n167) );
  N1M1P U41 ( .A(Packet_In[13]), .Z(n173) );
  N1M1P U42 ( .A(Packet_In[14]), .Z(n175) );
  N1M1P U43 ( .A(Packet_In[3]), .Z(n153) );
  N1M1P U44 ( .A(Packet_In[9]), .Z(n165) );
  N1M1P U45 ( .A(Packet_In[11]), .Z(n169) );
  N1M1P U46 ( .A(Packet_In[19]), .Z(n185) );
  N1M1P U47 ( .A(Packet_In[5]), .Z(n157) );
  N1M1P U48 ( .A(Packet_In[4]), .Z(n155) );
  N1M1P U49 ( .A(Packet_In[7]), .Z(n161) );
  N1M1P U50 ( .A(Packet_In[30]), .Z(n207) );
  N1M1P U51 ( .A(Packet_In[0]), .Z(n147) );
  N1M1P U52 ( .A(Packet_In[2]), .Z(n151) );
  N1M1P U53 ( .A(Packet_In[16]), .Z(n179) );
  N1M1P U54 ( .A(Packet_In[8]), .Z(n163) );
  N1M1P U55 ( .A(Packet_In[18]), .Z(n183) );
  N1M1P U56 ( .A(Packet_In[1]), .Z(n149) );
  N1M1P U57 ( .A(Packet_In[6]), .Z(n159) );
  N1M1P U58 ( .A(Packet_In[17]), .Z(n181) );
  N1M1P U59 ( .A(Packet_In[15]), .Z(n177) );
  BUFM2P U60 ( .A(n100), .Z(n11) );
  BUFM2P U61 ( .A(n60), .Z(n7) );
  BUFM2P U62 ( .A(n136), .Z(n13) );
  BUFM2P U63 ( .A(n136), .Z(n12) );
  BUFM2P U64 ( .A(n373), .Z(n14) );
  BUFM2P U65 ( .A(n373), .Z(n15) );
  BUFM2P U66 ( .A(n59), .Z(n6) );
  BUFM2P U67 ( .A(n59), .Z(n5) );
  BUFM2P U68 ( .A(n59), .Z(n4) );
  N1M2P U69 ( .A(n21), .Z(n142) );
  BUFM2P U70 ( .A(n97), .Z(n9) );
  BUFM2P U71 ( .A(n97), .Z(n8) );
  N1M2P U72 ( .A(n65), .Z(n97) );
  OAI211M1P U73 ( .A(n379), .B(n140), .C(n3), .D(n65), .Z(n100) );
  NR2M1P U74 ( .A(n140), .B(n3), .Z(n378) );
  NR2M1P U75 ( .A(n21), .B(n378), .Z(n377) );
  AOI22CDNM1P U76 ( .A(n377), .B(n26), .C(n377), .D(n26), .Z(n372) );
  N1M1P U77 ( .A(n378), .Z(n20) );
  AOI22M1P U78 ( .A(Count[0]), .B(n142), .C(n20), .D(n26), .Z(n17) );
  AOI22CDNM1P U79 ( .A(Count[1]), .B(n17), .C(n17), .D(Count[1]), .Z(n371) );
  ND3M1P U80 ( .A(n26), .B(n22), .C(n25), .Z(n63) );
  ND2M1P U81 ( .A(Count[1]), .B(Read_Ack), .Z(n16) );
  OAI211M1P U82 ( .A(Count[1]), .B(n142), .C(n17), .D(n16), .Z(n18) );
  AOI22M1P U83 ( .A(n21), .B(n143), .C(Count[2]), .D(n18), .Z(n19) );
  OAI21M1P U84 ( .A(n63), .B(n20), .C(n19), .Z(n370) );
  AOI22CDNM1P U85 ( .A(n23), .B(n376), .C(\Queue[4][31] ), .D(n23), .Z(n369)
         );
  AOI22CDNM1P U86 ( .A(n23), .B(n147), .C(\Queue[4][0] ), .D(n23), .Z(n368) );
  AOI22CDNM1P U87 ( .A(n23), .B(n149), .C(\Queue[4][1] ), .D(n23), .Z(n367) );
  AOI22CDNM1P U88 ( .A(n23), .B(n151), .C(\Queue[4][2] ), .D(n23), .Z(n366) );
  AOI22CDNM1P U89 ( .A(n23), .B(n153), .C(\Queue[4][3] ), .D(n23), .Z(n365) );
  AOI22CDNM1P U90 ( .A(n23), .B(n155), .C(\Queue[4][4] ), .D(n23), .Z(n364) );
  AOI22CDNM1P U91 ( .A(n23), .B(n157), .C(\Queue[4][5] ), .D(n23), .Z(n363) );
  AOI22CDNM1P U92 ( .A(n23), .B(n159), .C(\Queue[4][6] ), .D(n23), .Z(n362) );
  AOI22CDNM1P U93 ( .A(n23), .B(n161), .C(\Queue[4][7] ), .D(n23), .Z(n361) );
  AOI22CDNM1P U94 ( .A(n23), .B(n163), .C(\Queue[4][8] ), .D(n23), .Z(n360) );
  AOI22CDNM1P U95 ( .A(n23), .B(n165), .C(\Queue[4][9] ), .D(n23), .Z(n359) );
  AOI22CDNM1P U96 ( .A(n23), .B(n167), .C(\Queue[4][10] ), .D(n23), .Z(n358)
         );
  AOI22CDNM1P U97 ( .A(n23), .B(n169), .C(\Queue[4][11] ), .D(n23), .Z(n357)
         );
  AOI22CDNM1P U98 ( .A(n23), .B(n171), .C(\Queue[4][12] ), .D(n23), .Z(n356)
         );
  AOI22CDNM1P U99 ( .A(n23), .B(n173), .C(\Queue[4][13] ), .D(n23), .Z(n355)
         );
  AOI22CDNM1P U100 ( .A(n23), .B(n175), .C(\Queue[4][14] ), .D(n23), .Z(n354)
         );
  AOI22CDNM1P U101 ( .A(n23), .B(n177), .C(\Queue[4][15] ), .D(n23), .Z(n353)
         );
  AOI22CDNM1P U102 ( .A(n23), .B(n179), .C(\Queue[4][16] ), .D(n23), .Z(n352)
         );
  AOI22CDNM1P U103 ( .A(n23), .B(n181), .C(\Queue[4][17] ), .D(n23), .Z(n351)
         );
  AOI22CDNM1P U104 ( .A(n23), .B(n183), .C(\Queue[4][18] ), .D(n23), .Z(n350)
         );
  AOI22CDNM1P U105 ( .A(n23), .B(n185), .C(\Queue[4][19] ), .D(n23), .Z(n349)
         );
  AOI22CDNM1P U106 ( .A(n23), .B(n187), .C(\Queue[4][20] ), .D(n23), .Z(n348)
         );
  AOI22CDNM1P U107 ( .A(n23), .B(n189), .C(\Queue[4][21] ), .D(n23), .Z(n347)
         );
  AOI22CDNM1P U108 ( .A(n23), .B(n191), .C(\Queue[4][22] ), .D(n23), .Z(n346)
         );
  AOI22CDNM1P U109 ( .A(n23), .B(n193), .C(\Queue[4][23] ), .D(n23), .Z(n345)
         );
  AOI22CDNM1P U110 ( .A(n23), .B(n195), .C(\Queue[4][24] ), .D(n23), .Z(n344)
         );
  AOI22CDNM1P U111 ( .A(n23), .B(n197), .C(\Queue[4][25] ), .D(n23), .Z(n343)
         );
  AOI22CDNM1P U112 ( .A(n23), .B(n199), .C(\Queue[4][26] ), .D(n23), .Z(n342)
         );
  AOI22CDNM1P U113 ( .A(n23), .B(n201), .C(\Queue[4][27] ), .D(n23), .Z(n341)
         );
  AOI22CDNM1P U114 ( .A(n23), .B(n203), .C(\Queue[4][28] ), .D(n23), .Z(n340)
         );
  AOI22CDNM1P U115 ( .A(n23), .B(n205), .C(\Queue[4][29] ), .D(n23), .Z(n339)
         );
  AOI22CDNM1P U116 ( .A(n23), .B(n207), .C(\Queue[4][30] ), .D(n23), .Z(n338)
         );
  OAI22CDNM1P U117 ( .A(n142), .B(n24), .C(n377), .D(Full), .Z(n337) );
  OA21M1P U118 ( .A(n142), .B(n379), .C(Rst_n), .Z(n27) );
  OAI21M1P U119 ( .A(n3), .B(Read_Ack), .C(n27), .Z(n59) );
  AOI22M1P U120 ( .A(\Queue[2][0] ), .B(n60), .C(\Queue[1][0] ), .D(n4), .Z(
        n28) );
  OAI21M1P U121 ( .A(n147), .B(n62), .C(n28), .Z(n336) );
  AOI22M1P U122 ( .A(n7), .B(\Queue[2][1] ), .C(\Queue[1][1] ), .D(n4), .Z(n29) );
  OAI21M1P U123 ( .A(n62), .B(n149), .C(n29), .Z(n335) );
  AOI22M1P U124 ( .A(n60), .B(\Queue[2][2] ), .C(\Queue[1][2] ), .D(n4), .Z(
        n30) );
  OAI21M1P U125 ( .A(n62), .B(n151), .C(n30), .Z(n334) );
  AOI22M1P U126 ( .A(n60), .B(\Queue[2][3] ), .C(\Queue[1][3] ), .D(n4), .Z(
        n31) );
  OAI21M1P U127 ( .A(n62), .B(n153), .C(n31), .Z(n333) );
  AOI22M1P U128 ( .A(n60), .B(\Queue[2][4] ), .C(\Queue[1][4] ), .D(n4), .Z(
        n32) );
  OAI21M1P U129 ( .A(n62), .B(n155), .C(n32), .Z(n332) );
  AOI22M1P U130 ( .A(n60), .B(\Queue[2][5] ), .C(\Queue[1][5] ), .D(n4), .Z(
        n33) );
  OAI21M1P U131 ( .A(n62), .B(n157), .C(n33), .Z(n331) );
  AOI22M1P U132 ( .A(n60), .B(\Queue[2][6] ), .C(\Queue[1][6] ), .D(n4), .Z(
        n34) );
  OAI21M1P U133 ( .A(n62), .B(n159), .C(n34), .Z(n330) );
  AOI22M1P U134 ( .A(n60), .B(\Queue[2][7] ), .C(\Queue[1][7] ), .D(n4), .Z(
        n35) );
  OAI21M1P U135 ( .A(n62), .B(n161), .C(n35), .Z(n329) );
  AOI22M1P U136 ( .A(n60), .B(\Queue[2][8] ), .C(\Queue[1][8] ), .D(n4), .Z(
        n36) );
  OAI21M1P U137 ( .A(n62), .B(n163), .C(n36), .Z(n328) );
  AOI22M1P U138 ( .A(n60), .B(\Queue[2][9] ), .C(\Queue[1][9] ), .D(n5), .Z(
        n37) );
  OAI21M1P U139 ( .A(n62), .B(n165), .C(n37), .Z(n327) );
  AOI22M1P U140 ( .A(n60), .B(\Queue[2][10] ), .C(\Queue[1][10] ), .D(n5), .Z(
        n38) );
  OAI21M1P U141 ( .A(n62), .B(n167), .C(n38), .Z(n326) );
  AOI22M1P U142 ( .A(n60), .B(\Queue[2][11] ), .C(\Queue[1][11] ), .D(n5), .Z(
        n39) );
  OAI21M1P U143 ( .A(n62), .B(n169), .C(n39), .Z(n325) );
  AOI22M1P U144 ( .A(n7), .B(\Queue[2][12] ), .C(\Queue[1][12] ), .D(n5), .Z(
        n40) );
  OAI21M1P U145 ( .A(n62), .B(n171), .C(n40), .Z(n324) );
  AOI22M1P U146 ( .A(n7), .B(\Queue[2][13] ), .C(\Queue[1][13] ), .D(n5), .Z(
        n41) );
  OAI21M1P U147 ( .A(n62), .B(n173), .C(n41), .Z(n323) );
  AOI22M1P U148 ( .A(n7), .B(\Queue[2][14] ), .C(\Queue[1][14] ), .D(n5), .Z(
        n42) );
  OAI21M1P U149 ( .A(n62), .B(n175), .C(n42), .Z(n322) );
  AOI22M1P U150 ( .A(n7), .B(\Queue[2][15] ), .C(\Queue[1][15] ), .D(n5), .Z(
        n43) );
  OAI21M1P U151 ( .A(n62), .B(n177), .C(n43), .Z(n321) );
  AOI22M1P U152 ( .A(n7), .B(\Queue[2][16] ), .C(\Queue[1][16] ), .D(n5), .Z(
        n44) );
  OAI21M1P U153 ( .A(n62), .B(n179), .C(n44), .Z(n320) );
  AOI22M1P U154 ( .A(n7), .B(\Queue[2][17] ), .C(\Queue[1][17] ), .D(n5), .Z(
        n45) );
  OAI21M1P U155 ( .A(n62), .B(n181), .C(n45), .Z(n319) );
  AOI22M1P U156 ( .A(n7), .B(\Queue[2][18] ), .C(\Queue[1][18] ), .D(n6), .Z(
        n46) );
  OAI21M1P U157 ( .A(n62), .B(n183), .C(n46), .Z(n318) );
  AOI22M1P U158 ( .A(n7), .B(\Queue[2][19] ), .C(\Queue[1][19] ), .D(n6), .Z(
        n47) );
  OAI21M1P U159 ( .A(n62), .B(n185), .C(n47), .Z(n317) );
  AOI22M1P U160 ( .A(n7), .B(\Queue[2][20] ), .C(\Queue[1][20] ), .D(n6), .Z(
        n48) );
  OAI21M1P U161 ( .A(n62), .B(n187), .C(n48), .Z(n316) );
  AOI22M1P U162 ( .A(n7), .B(\Queue[2][21] ), .C(\Queue[1][21] ), .D(n6), .Z(
        n49) );
  OAI21M1P U163 ( .A(n62), .B(n189), .C(n49), .Z(n315) );
  AOI22M1P U164 ( .A(n7), .B(\Queue[2][22] ), .C(\Queue[1][22] ), .D(n6), .Z(
        n50) );
  OAI21M1P U165 ( .A(n62), .B(n191), .C(n50), .Z(n314) );
  AOI22M1P U166 ( .A(n7), .B(\Queue[2][23] ), .C(\Queue[1][23] ), .D(n6), .Z(
        n51) );
  OAI21M1P U167 ( .A(n62), .B(n193), .C(n51), .Z(n313) );
  AOI22M1P U168 ( .A(n60), .B(\Queue[2][24] ), .C(\Queue[1][24] ), .D(n6), .Z(
        n52) );
  OAI21M1P U169 ( .A(n62), .B(n195), .C(n52), .Z(n312) );
  AOI22M1P U170 ( .A(n60), .B(\Queue[2][25] ), .C(\Queue[1][25] ), .D(n6), .Z(
        n53) );
  OAI21M1P U171 ( .A(n62), .B(n197), .C(n53), .Z(n311) );
  AOI22M1P U172 ( .A(n60), .B(\Queue[2][26] ), .C(\Queue[1][26] ), .D(n6), .Z(
        n54) );
  OAI21M1P U173 ( .A(n62), .B(n199), .C(n54), .Z(n310) );
  AOI22M1P U174 ( .A(n60), .B(\Queue[2][27] ), .C(\Queue[1][27] ), .D(n6), .Z(
        n55) );
  OAI21M1P U175 ( .A(n62), .B(n201), .C(n55), .Z(n309) );
  AOI22M1P U176 ( .A(n60), .B(\Queue[2][28] ), .C(\Queue[1][28] ), .D(n4), .Z(
        n56) );
  OAI21M1P U177 ( .A(n62), .B(n203), .C(n56), .Z(n308) );
  AOI22M1P U178 ( .A(n60), .B(\Queue[2][29] ), .C(\Queue[1][29] ), .D(n5), .Z(
        n57) );
  OAI21M1P U179 ( .A(n62), .B(n205), .C(n57), .Z(n307) );
  AOI22M1P U180 ( .A(n60), .B(\Queue[2][30] ), .C(\Queue[1][30] ), .D(n6), .Z(
        n58) );
  OAI21M1P U181 ( .A(n62), .B(n207), .C(n58), .Z(n306) );
  AOI22M1P U182 ( .A(n60), .B(\Queue[2][31] ), .C(\Queue[1][31] ), .D(n4), .Z(
        n61) );
  OAI21M1P U183 ( .A(n62), .B(n376), .C(n61), .Z(n305) );
  OAI21M1P U184 ( .A(n64), .B(n63), .C(n144), .Z(n65) );
  AOI22M1P U185 ( .A(\Queue[1][0] ), .B(n98), .C(n8), .D(Packet_Out[0]), .Z(
        n66) );
  OAI21M1P U186 ( .A(n147), .B(n10), .C(n66), .Z(n304) );
  AOI22M1P U187 ( .A(\Queue[1][1] ), .B(n98), .C(n8), .D(Packet_Out[1]), .Z(
        n67) );
  OAI21M1P U188 ( .A(n149), .B(n10), .C(n67), .Z(n303) );
  AOI22M1P U189 ( .A(\Queue[1][2] ), .B(n98), .C(n8), .D(Packet_Out[2]), .Z(
        n68) );
  OAI21M1P U190 ( .A(n151), .B(n10), .C(n68), .Z(n302) );
  AOI22M1P U191 ( .A(\Queue[1][3] ), .B(n98), .C(n8), .D(Packet_Out[3]), .Z(
        n69) );
  OAI21M1P U192 ( .A(n153), .B(n10), .C(n69), .Z(n301) );
  AOI22M1P U193 ( .A(\Queue[1][4] ), .B(n98), .C(n8), .D(Packet_Out[4]), .Z(
        n70) );
  OAI21M1P U194 ( .A(n155), .B(n10), .C(n70), .Z(n300) );
  AOI22M1P U195 ( .A(\Queue[1][5] ), .B(n98), .C(n8), .D(Packet_Out[5]), .Z(
        n71) );
  OAI21M1P U196 ( .A(n157), .B(n10), .C(n71), .Z(n299) );
  AOI22M1P U197 ( .A(\Queue[1][6] ), .B(n98), .C(n8), .D(Packet_Out[6]), .Z(
        n72) );
  OAI21M1P U198 ( .A(n159), .B(n10), .C(n72), .Z(n298) );
  AOI22M1P U199 ( .A(\Queue[1][7] ), .B(n98), .C(n8), .D(Packet_Out[7]), .Z(
        n73) );
  OAI21M1P U200 ( .A(n161), .B(n10), .C(n73), .Z(n297) );
  AOI22M1P U201 ( .A(\Queue[1][8] ), .B(n98), .C(n8), .D(Packet_Out[8]), .Z(
        n74) );
  OAI21M1P U202 ( .A(n163), .B(n10), .C(n74), .Z(n296) );
  AOI22M1P U203 ( .A(\Queue[1][9] ), .B(n98), .C(n8), .D(Packet_Out[9]), .Z(
        n75) );
  OAI21M1P U204 ( .A(n165), .B(n10), .C(n75), .Z(n295) );
  AOI22M1P U205 ( .A(\Queue[1][10] ), .B(n98), .C(n97), .D(Packet_Out[10]), 
        .Z(n76) );
  OAI21M1P U206 ( .A(n167), .B(n10), .C(n76), .Z(n294) );
  AOI22M1P U207 ( .A(\Queue[1][11] ), .B(n98), .C(n97), .D(Packet_Out[11]), 
        .Z(n77) );
  OAI21M1P U208 ( .A(n169), .B(n10), .C(n77), .Z(n293) );
  AOI22M1P U209 ( .A(\Queue[1][12] ), .B(n98), .C(n97), .D(Packet_Out[12]), 
        .Z(n78) );
  OAI21M1P U210 ( .A(n171), .B(n10), .C(n78), .Z(n292) );
  AOI22M1P U211 ( .A(\Queue[1][13] ), .B(n98), .C(n97), .D(Packet_Out[13]), 
        .Z(n79) );
  OAI21M1P U212 ( .A(n173), .B(n10), .C(n79), .Z(n291) );
  AOI22M1P U213 ( .A(\Queue[1][14] ), .B(n98), .C(n97), .D(Packet_Out[14]), 
        .Z(n80) );
  OAI21M1P U214 ( .A(n175), .B(n10), .C(n80), .Z(n290) );
  AOI22M1P U215 ( .A(\Queue[1][15] ), .B(n98), .C(n97), .D(Packet_Out[15]), 
        .Z(n81) );
  OAI21M1P U216 ( .A(n177), .B(n10), .C(n81), .Z(n289) );
  AOI22M1P U217 ( .A(\Queue[1][16] ), .B(n98), .C(n97), .D(Packet_Out[16]), 
        .Z(n82) );
  OAI21M1P U218 ( .A(n179), .B(n10), .C(n82), .Z(n288) );
  AOI22M1P U219 ( .A(\Queue[1][17] ), .B(n98), .C(n97), .D(Packet_Out[17]), 
        .Z(n83) );
  OAI21M1P U220 ( .A(n181), .B(n10), .C(n83), .Z(n287) );
  AOI22M1P U221 ( .A(\Queue[1][18] ), .B(n98), .C(n97), .D(Packet_Out[18]), 
        .Z(n84) );
  OAI21M1P U222 ( .A(n183), .B(n10), .C(n84), .Z(n286) );
  AOI22M1P U223 ( .A(\Queue[1][19] ), .B(n98), .C(n97), .D(Packet_Out[19]), 
        .Z(n85) );
  OAI21M1P U224 ( .A(n185), .B(n10), .C(n85), .Z(n285) );
  AOI22M1P U225 ( .A(\Queue[1][20] ), .B(n98), .C(n9), .D(Packet_Out[20]), .Z(
        n86) );
  OAI21M1P U226 ( .A(n187), .B(n11), .C(n86), .Z(n284) );
  AOI22M1P U227 ( .A(\Queue[1][21] ), .B(n98), .C(n9), .D(Packet_Out[21]), .Z(
        n87) );
  OAI21M1P U228 ( .A(n189), .B(n11), .C(n87), .Z(n283) );
  AOI22M1P U229 ( .A(\Queue[1][22] ), .B(n98), .C(n9), .D(Packet_Out[22]), .Z(
        n88) );
  OAI21M1P U230 ( .A(n191), .B(n11), .C(n88), .Z(n282) );
  AOI22M1P U231 ( .A(\Queue[1][23] ), .B(n98), .C(n9), .D(Packet_Out[23]), .Z(
        n89) );
  OAI21M1P U232 ( .A(n193), .B(n11), .C(n89), .Z(n281) );
  AOI22M1P U233 ( .A(\Queue[1][24] ), .B(n98), .C(n9), .D(Packet_Out[24]), .Z(
        n90) );
  OAI21M1P U234 ( .A(n195), .B(n11), .C(n90), .Z(n280) );
  AOI22M1P U235 ( .A(\Queue[1][25] ), .B(n98), .C(n9), .D(Packet_Out[25]), .Z(
        n91) );
  OAI21M1P U236 ( .A(n197), .B(n11), .C(n91), .Z(n279) );
  AOI22M1P U237 ( .A(\Queue[1][26] ), .B(n98), .C(n9), .D(Packet_Out[26]), .Z(
        n92) );
  OAI21M1P U238 ( .A(n199), .B(n11), .C(n92), .Z(n278) );
  AOI22M1P U239 ( .A(\Queue[1][27] ), .B(n98), .C(n9), .D(Packet_Out[27]), .Z(
        n93) );
  OAI21M1P U240 ( .A(n201), .B(n11), .C(n93), .Z(n277) );
  AOI22M1P U241 ( .A(\Queue[1][28] ), .B(n98), .C(n9), .D(Packet_Out[28]), .Z(
        n94) );
  OAI21M1P U242 ( .A(n203), .B(n11), .C(n94), .Z(n276) );
  AOI22M1P U243 ( .A(\Queue[1][29] ), .B(n98), .C(n9), .D(Packet_Out[29]), .Z(
        n95) );
  OAI21M1P U244 ( .A(n205), .B(n11), .C(n95), .Z(n275) );
  AOI22M1P U245 ( .A(\Queue[1][30] ), .B(n98), .C(n9), .D(Packet_Out[30]), .Z(
        n96) );
  OAI21M1P U246 ( .A(n207), .B(n10), .C(n96), .Z(n274) );
  AOI22M1P U247 ( .A(\Queue[1][31] ), .B(n98), .C(n8), .D(Packet_Out[31]), .Z(
        n99) );
  OAI21M1P U248 ( .A(n376), .B(n11), .C(n99), .Z(n273) );
  OA21M1P U249 ( .A(n142), .B(n103), .C(Rst_n), .Z(n101) );
  ND2M1P U250 ( .A(n102), .B(n140), .Z(n141) );
  AOI22M1P U251 ( .A(\Queue[2][0] ), .B(n136), .C(\Queue[3][0] ), .D(n135), 
        .Z(n104) );
  OAI21M1P U252 ( .A(n147), .B(n138), .C(n104), .Z(n272) );
  AOI22M1P U253 ( .A(\Queue[2][1] ), .B(n136), .C(n135), .D(\Queue[3][1] ), 
        .Z(n105) );
  OAI21M1P U254 ( .A(n149), .B(n138), .C(n105), .Z(n271) );
  AOI22M1P U255 ( .A(\Queue[2][2] ), .B(n136), .C(n135), .D(\Queue[3][2] ), 
        .Z(n106) );
  OAI21M1P U256 ( .A(n151), .B(n138), .C(n106), .Z(n270) );
  AOI22M1P U257 ( .A(\Queue[2][3] ), .B(n136), .C(n135), .D(\Queue[3][3] ), 
        .Z(n107) );
  OAI21M1P U258 ( .A(n153), .B(n138), .C(n107), .Z(n269) );
  AOI22M1P U259 ( .A(\Queue[2][4] ), .B(n136), .C(n135), .D(\Queue[3][4] ), 
        .Z(n108) );
  OAI21M1P U260 ( .A(n155), .B(n138), .C(n108), .Z(n268) );
  AOI22M1P U261 ( .A(\Queue[2][5] ), .B(n136), .C(n135), .D(\Queue[3][5] ), 
        .Z(n109) );
  OAI21M1P U262 ( .A(n157), .B(n138), .C(n109), .Z(n267) );
  AOI22M1P U263 ( .A(\Queue[2][6] ), .B(n12), .C(n135), .D(\Queue[3][6] ), .Z(
        n110) );
  OAI21M1P U264 ( .A(n159), .B(n138), .C(n110), .Z(n266) );
  AOI22M1P U265 ( .A(\Queue[2][7] ), .B(n13), .C(n135), .D(\Queue[3][7] ), .Z(
        n111) );
  OAI21M1P U266 ( .A(n161), .B(n138), .C(n111), .Z(n265) );
  AOI22M1P U267 ( .A(\Queue[2][8] ), .B(n12), .C(n135), .D(\Queue[3][8] ), .Z(
        n112) );
  OAI21M1P U268 ( .A(n163), .B(n138), .C(n112), .Z(n264) );
  AOI22M1P U269 ( .A(\Queue[2][9] ), .B(n13), .C(n135), .D(\Queue[3][9] ), .Z(
        n113) );
  OAI21M1P U270 ( .A(n165), .B(n138), .C(n113), .Z(n263) );
  AOI22M1P U271 ( .A(\Queue[2][10] ), .B(n12), .C(n135), .D(\Queue[3][10] ), 
        .Z(n114) );
  OAI21M1P U272 ( .A(n167), .B(n138), .C(n114), .Z(n262) );
  AOI22M1P U273 ( .A(\Queue[2][11] ), .B(n12), .C(n135), .D(\Queue[3][11] ), 
        .Z(n115) );
  OAI21M1P U274 ( .A(n169), .B(n138), .C(n115), .Z(n261) );
  AOI22M1P U275 ( .A(\Queue[2][12] ), .B(n12), .C(n135), .D(\Queue[3][12] ), 
        .Z(n116) );
  OAI21M1P U276 ( .A(n171), .B(n138), .C(n116), .Z(n260) );
  AOI22M1P U277 ( .A(\Queue[2][13] ), .B(n12), .C(n135), .D(\Queue[3][13] ), 
        .Z(n117) );
  OAI21M1P U278 ( .A(n173), .B(n138), .C(n117), .Z(n259) );
  AOI22M1P U279 ( .A(\Queue[2][14] ), .B(n12), .C(n135), .D(\Queue[3][14] ), 
        .Z(n118) );
  OAI21M1P U280 ( .A(n175), .B(n138), .C(n118), .Z(n258) );
  AOI22M1P U281 ( .A(\Queue[2][15] ), .B(n12), .C(n135), .D(\Queue[3][15] ), 
        .Z(n119) );
  OAI21M1P U282 ( .A(n177), .B(n138), .C(n119), .Z(n257) );
  AOI22M1P U283 ( .A(\Queue[2][16] ), .B(n12), .C(n135), .D(\Queue[3][16] ), 
        .Z(n120) );
  OAI21M1P U284 ( .A(n179), .B(n138), .C(n120), .Z(n256) );
  AOI22M1P U285 ( .A(\Queue[2][17] ), .B(n12), .C(n135), .D(\Queue[3][17] ), 
        .Z(n121) );
  OAI21M1P U286 ( .A(n181), .B(n138), .C(n121), .Z(n255) );
  AOI22M1P U287 ( .A(\Queue[2][18] ), .B(n12), .C(n135), .D(\Queue[3][18] ), 
        .Z(n122) );
  OAI21M1P U288 ( .A(n183), .B(n138), .C(n122), .Z(n254) );
  AOI22M1P U289 ( .A(\Queue[2][19] ), .B(n12), .C(n135), .D(\Queue[3][19] ), 
        .Z(n123) );
  OAI21M1P U290 ( .A(n185), .B(n138), .C(n123), .Z(n253) );
  AOI22M1P U291 ( .A(\Queue[2][20] ), .B(n13), .C(n135), .D(\Queue[3][20] ), 
        .Z(n124) );
  OAI21M1P U292 ( .A(n187), .B(n138), .C(n124), .Z(n252) );
  AOI22M1P U293 ( .A(\Queue[2][21] ), .B(n13), .C(n135), .D(\Queue[3][21] ), 
        .Z(n125) );
  OAI21M1P U294 ( .A(n189), .B(n138), .C(n125), .Z(n251) );
  AOI22M1P U295 ( .A(\Queue[2][22] ), .B(n13), .C(n135), .D(\Queue[3][22] ), 
        .Z(n126) );
  OAI21M1P U296 ( .A(n191), .B(n138), .C(n126), .Z(n250) );
  AOI22M1P U297 ( .A(\Queue[2][23] ), .B(n13), .C(n135), .D(\Queue[3][23] ), 
        .Z(n127) );
  OAI21M1P U298 ( .A(n193), .B(n138), .C(n127), .Z(n249) );
  AOI22M1P U299 ( .A(\Queue[2][24] ), .B(n13), .C(n135), .D(\Queue[3][24] ), 
        .Z(n128) );
  OAI21M1P U300 ( .A(n195), .B(n138), .C(n128), .Z(n248) );
  AOI22M1P U301 ( .A(\Queue[2][25] ), .B(n13), .C(n135), .D(\Queue[3][25] ), 
        .Z(n129) );
  OAI21M1P U302 ( .A(n197), .B(n138), .C(n129), .Z(n247) );
  AOI22M1P U303 ( .A(\Queue[2][26] ), .B(n13), .C(n135), .D(\Queue[3][26] ), 
        .Z(n130) );
  OAI21M1P U304 ( .A(n199), .B(n138), .C(n130), .Z(n246) );
  AOI22M1P U305 ( .A(\Queue[2][27] ), .B(n13), .C(n135), .D(\Queue[3][27] ), 
        .Z(n131) );
  OAI21M1P U306 ( .A(n201), .B(n138), .C(n131), .Z(n245) );
  AOI22M1P U307 ( .A(\Queue[2][28] ), .B(n13), .C(n135), .D(\Queue[3][28] ), 
        .Z(n132) );
  OAI21M1P U308 ( .A(n203), .B(n138), .C(n132), .Z(n244) );
  AOI22M1P U309 ( .A(\Queue[2][29] ), .B(n13), .C(n135), .D(\Queue[3][29] ), 
        .Z(n133) );
  OAI21M1P U310 ( .A(n205), .B(n138), .C(n133), .Z(n243) );
  AOI22M1P U311 ( .A(\Queue[2][30] ), .B(n12), .C(n135), .D(\Queue[3][30] ), 
        .Z(n134) );
  OAI21M1P U312 ( .A(n207), .B(n138), .C(n134), .Z(n242) );
  AOI22M1P U313 ( .A(\Queue[2][31] ), .B(n13), .C(n135), .D(\Queue[3][31] ), 
        .Z(n137) );
  OAI21M1P U314 ( .A(n376), .B(n138), .C(n137), .Z(n241) );
  OA21M1P U315 ( .A(n142), .B(n143), .C(Rst_n), .Z(n139) );
  AOI22M1P U316 ( .A(\Queue[3][0] ), .B(n15), .C(n208), .D(\Queue[4][0] ), .Z(
        n146) );
  OAI21M1P U317 ( .A(n147), .B(n375), .C(n146), .Z(n240) );
  AOI22M1P U318 ( .A(\Queue[3][1] ), .B(n373), .C(n208), .D(\Queue[4][1] ), 
        .Z(n148) );
  OAI21M1P U319 ( .A(n149), .B(n375), .C(n148), .Z(n239) );
  AOI22M1P U320 ( .A(\Queue[3][2] ), .B(n373), .C(n208), .D(\Queue[4][2] ), 
        .Z(n150) );
  OAI21M1P U321 ( .A(n151), .B(n375), .C(n150), .Z(n238) );
  AOI22M1P U322 ( .A(\Queue[3][3] ), .B(n373), .C(n208), .D(\Queue[4][3] ), 
        .Z(n152) );
  OAI21M1P U323 ( .A(n153), .B(n375), .C(n152), .Z(n237) );
  AOI22M1P U324 ( .A(\Queue[3][4] ), .B(n373), .C(n208), .D(\Queue[4][4] ), 
        .Z(n154) );
  OAI21M1P U325 ( .A(n155), .B(n375), .C(n154), .Z(n236) );
  AOI22M1P U326 ( .A(\Queue[3][5] ), .B(n373), .C(n208), .D(\Queue[4][5] ), 
        .Z(n156) );
  OAI21M1P U327 ( .A(n157), .B(n375), .C(n156), .Z(n235) );
  AOI22M1P U328 ( .A(\Queue[3][6] ), .B(n373), .C(n208), .D(\Queue[4][6] ), 
        .Z(n158) );
  OAI21M1P U329 ( .A(n159), .B(n375), .C(n158), .Z(n234) );
  AOI22M1P U330 ( .A(\Queue[3][7] ), .B(n14), .C(n208), .D(\Queue[4][7] ), .Z(
        n160) );
  OAI21M1P U331 ( .A(n161), .B(n375), .C(n160), .Z(n233) );
  AOI22M1P U332 ( .A(\Queue[3][8] ), .B(n15), .C(n208), .D(\Queue[4][8] ), .Z(
        n162) );
  OAI21M1P U333 ( .A(n163), .B(n375), .C(n162), .Z(n232) );
  AOI22M1P U334 ( .A(\Queue[3][9] ), .B(n14), .C(n208), .D(\Queue[4][9] ), .Z(
        n164) );
  OAI21M1P U335 ( .A(n165), .B(n375), .C(n164), .Z(n231) );
  AOI22M1P U336 ( .A(\Queue[3][10] ), .B(n14), .C(n208), .D(\Queue[4][10] ), 
        .Z(n166) );
  OAI21M1P U337 ( .A(n167), .B(n375), .C(n166), .Z(n230) );
  AOI22M1P U338 ( .A(\Queue[3][11] ), .B(n14), .C(n208), .D(\Queue[4][11] ), 
        .Z(n168) );
  OAI21M1P U339 ( .A(n169), .B(n375), .C(n168), .Z(n229) );
  AOI22M1P U340 ( .A(\Queue[3][12] ), .B(n14), .C(n208), .D(\Queue[4][12] ), 
        .Z(n170) );
  OAI21M1P U341 ( .A(n171), .B(n375), .C(n170), .Z(n228) );
  AOI22M1P U342 ( .A(\Queue[3][13] ), .B(n14), .C(n208), .D(\Queue[4][13] ), 
        .Z(n172) );
  OAI21M1P U343 ( .A(n173), .B(n375), .C(n172), .Z(n227) );
  AOI22M1P U344 ( .A(\Queue[3][14] ), .B(n14), .C(n208), .D(\Queue[4][14] ), 
        .Z(n174) );
  OAI21M1P U345 ( .A(n175), .B(n375), .C(n174), .Z(n226) );
  AOI22M1P U346 ( .A(\Queue[3][15] ), .B(n14), .C(n208), .D(\Queue[4][15] ), 
        .Z(n176) );
  OAI21M1P U347 ( .A(n177), .B(n375), .C(n176), .Z(n225) );
  AOI22M1P U348 ( .A(\Queue[3][16] ), .B(n14), .C(n208), .D(\Queue[4][16] ), 
        .Z(n178) );
  OAI21M1P U349 ( .A(n179), .B(n375), .C(n178), .Z(n224) );
  AOI22M1P U350 ( .A(\Queue[3][17] ), .B(n14), .C(n208), .D(\Queue[4][17] ), 
        .Z(n180) );
  OAI21M1P U351 ( .A(n181), .B(n375), .C(n180), .Z(n223) );
  AOI22M1P U352 ( .A(\Queue[3][18] ), .B(n14), .C(n208), .D(\Queue[4][18] ), 
        .Z(n182) );
  OAI21M1P U353 ( .A(n183), .B(n375), .C(n182), .Z(n222) );
  AOI22M1P U354 ( .A(\Queue[3][19] ), .B(n14), .C(n208), .D(\Queue[4][19] ), 
        .Z(n184) );
  OAI21M1P U355 ( .A(n185), .B(n375), .C(n184), .Z(n221) );
  AOI22M1P U356 ( .A(\Queue[3][20] ), .B(n15), .C(n208), .D(\Queue[4][20] ), 
        .Z(n186) );
  OAI21M1P U357 ( .A(n187), .B(n375), .C(n186), .Z(n220) );
  AOI22M1P U358 ( .A(\Queue[3][21] ), .B(n15), .C(n208), .D(\Queue[4][21] ), 
        .Z(n188) );
  OAI21M1P U359 ( .A(n189), .B(n375), .C(n188), .Z(n219) );
  AOI22M1P U360 ( .A(\Queue[3][22] ), .B(n15), .C(n208), .D(\Queue[4][22] ), 
        .Z(n190) );
  OAI21M1P U361 ( .A(n191), .B(n375), .C(n190), .Z(n218) );
  AOI22M1P U362 ( .A(\Queue[3][23] ), .B(n15), .C(n208), .D(\Queue[4][23] ), 
        .Z(n192) );
  OAI21M1P U363 ( .A(n193), .B(n375), .C(n192), .Z(n217) );
  AOI22M1P U364 ( .A(\Queue[3][24] ), .B(n15), .C(n208), .D(\Queue[4][24] ), 
        .Z(n194) );
  OAI21M1P U365 ( .A(n195), .B(n375), .C(n194), .Z(n216) );
  AOI22M1P U366 ( .A(\Queue[3][25] ), .B(n15), .C(n208), .D(\Queue[4][25] ), 
        .Z(n196) );
  OAI21M1P U367 ( .A(n197), .B(n375), .C(n196), .Z(n215) );
  AOI22M1P U368 ( .A(\Queue[3][26] ), .B(n15), .C(n208), .D(\Queue[4][26] ), 
        .Z(n198) );
  OAI21M1P U369 ( .A(n199), .B(n375), .C(n198), .Z(n214) );
  AOI22M1P U370 ( .A(\Queue[3][27] ), .B(n15), .C(n208), .D(\Queue[4][27] ), 
        .Z(n200) );
  OAI21M1P U371 ( .A(n201), .B(n375), .C(n200), .Z(n213) );
  AOI22M1P U372 ( .A(\Queue[3][28] ), .B(n15), .C(n208), .D(\Queue[4][28] ), 
        .Z(n202) );
  OAI21M1P U373 ( .A(n203), .B(n375), .C(n202), .Z(n212) );
  AOI22M1P U374 ( .A(\Queue[3][29] ), .B(n15), .C(n208), .D(\Queue[4][29] ), 
        .Z(n204) );
  OAI21M1P U375 ( .A(n205), .B(n375), .C(n204), .Z(n211) );
  AOI22M1P U376 ( .A(\Queue[3][30] ), .B(n14), .C(n208), .D(\Queue[4][30] ), 
        .Z(n206) );
  OAI21M1P U377 ( .A(n207), .B(n375), .C(n206), .Z(n210) );
  AOI22M1P U378 ( .A(\Queue[3][31] ), .B(n15), .C(n208), .D(\Queue[4][31] ), 
        .Z(n374) );
  OAI21M1P U379 ( .A(n376), .B(n375), .C(n374), .Z(n209) );
  N1M1P U380 ( .A(n2), .Z(Empty) );
  AOI22M1P U381 ( .A(n379), .B(n378), .C(n377), .D(Empty), .Z(n1) );
endmodule


module Packet_Queue_9 ( Clk_r, Rst_n, Packet_In, Read_Ack, Write_Ack, 
        Packet_Out, Empty, Full );
  input [31:0] Packet_In;
  output [31:0] Packet_Out;
  input Clk_r, Rst_n, Read_Ack, Write_Ack;
  output Empty, Full;
  wire   \Queue[4][31] , \Queue[4][30] , \Queue[4][29] , \Queue[4][28] ,
         \Queue[4][27] , \Queue[4][26] , \Queue[4][25] , \Queue[4][24] ,
         \Queue[4][23] , \Queue[4][22] , \Queue[4][21] , \Queue[4][20] ,
         \Queue[4][19] , \Queue[4][18] , \Queue[4][17] , \Queue[4][16] ,
         \Queue[4][15] , \Queue[4][14] , \Queue[4][13] , \Queue[4][12] ,
         \Queue[4][11] , \Queue[4][10] , \Queue[4][9] , \Queue[4][8] ,
         \Queue[4][7] , \Queue[4][6] , \Queue[4][5] , \Queue[4][4] ,
         \Queue[4][3] , \Queue[4][2] , \Queue[4][1] , \Queue[4][0] ,
         \Queue[3][31] , \Queue[3][30] , \Queue[3][29] , \Queue[3][28] ,
         \Queue[3][27] , \Queue[3][26] , \Queue[3][25] , \Queue[3][24] ,
         \Queue[3][23] , \Queue[3][22] , \Queue[3][21] , \Queue[3][20] ,
         \Queue[3][19] , \Queue[3][18] , \Queue[3][17] , \Queue[3][16] ,
         \Queue[3][15] , \Queue[3][14] , \Queue[3][13] , \Queue[3][12] ,
         \Queue[3][11] , \Queue[3][10] , \Queue[3][9] , \Queue[3][8] ,
         \Queue[3][7] , \Queue[3][6] , \Queue[3][5] , \Queue[3][4] ,
         \Queue[3][3] , \Queue[3][2] , \Queue[3][1] , \Queue[3][0] ,
         \Queue[2][31] , \Queue[2][30] , \Queue[2][29] , \Queue[2][28] ,
         \Queue[2][27] , \Queue[2][26] , \Queue[2][25] , \Queue[2][24] ,
         \Queue[2][23] , \Queue[2][22] , \Queue[2][21] , \Queue[2][20] ,
         \Queue[2][19] , \Queue[2][18] , \Queue[2][17] , \Queue[2][16] ,
         \Queue[2][15] , \Queue[2][14] , \Queue[2][13] , \Queue[2][12] ,
         \Queue[2][11] , \Queue[2][10] , \Queue[2][9] , \Queue[2][8] ,
         \Queue[2][7] , \Queue[2][6] , \Queue[2][5] , \Queue[2][4] ,
         \Queue[2][3] , \Queue[2][2] , \Queue[2][1] , \Queue[2][0] ,
         \Queue[1][31] , \Queue[1][30] , \Queue[1][29] , \Queue[1][28] ,
         \Queue[1][27] , \Queue[1][26] , \Queue[1][25] , \Queue[1][24] ,
         \Queue[1][23] , \Queue[1][22] , \Queue[1][21] , \Queue[1][20] ,
         \Queue[1][19] , \Queue[1][18] , \Queue[1][17] , \Queue[1][16] ,
         \Queue[1][15] , \Queue[1][14] , \Queue[1][13] , \Queue[1][12] ,
         \Queue[1][11] , \Queue[1][10] , \Queue[1][9] , \Queue[1][8] ,
         \Queue[1][7] , \Queue[1][6] , \Queue[1][5] , \Queue[1][4] ,
         \Queue[1][3] , \Queue[1][2] , \Queue[1][1] , \Queue[1][0] , n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539;
  wire   [2:0] Count;

  FDN2QM1P \Count_reg[0]  ( .D(n374), .CPN(Clk_r), .CD(Rst_n), .Q(Count[0]) );
  FDN2QM1P \Count_reg[1]  ( .D(n375), .CPN(Clk_r), .CD(Rst_n), .Q(Count[1]) );
  FDN2QM1P \Count_reg[2]  ( .D(n376), .CPN(Clk_r), .CD(Rst_n), .Q(Count[2]) );
  FDN1QM1P \Queue_reg[4][30]  ( .D(n408), .CPN(Clk_r), .Q(\Queue[4][30] ) );
  FDN1QM1P \Queue_reg[3][30]  ( .D(n536), .CPN(Clk_r), .Q(\Queue[3][30] ) );
  FDN1QM1P \Queue_reg[2][30]  ( .D(n504), .CPN(Clk_r), .Q(\Queue[2][30] ) );
  FDN1QM1P \Queue_reg[4][29]  ( .D(n407), .CPN(Clk_r), .Q(\Queue[4][29] ) );
  FDN1QM1P \Queue_reg[3][29]  ( .D(n535), .CPN(Clk_r), .Q(\Queue[3][29] ) );
  FDN1QM1P \Queue_reg[2][29]  ( .D(n503), .CPN(Clk_r), .Q(\Queue[2][29] ) );
  FDN1QM1P \Queue_reg[4][28]  ( .D(n406), .CPN(Clk_r), .Q(\Queue[4][28] ) );
  FDN1QM1P \Queue_reg[3][28]  ( .D(n534), .CPN(Clk_r), .Q(\Queue[3][28] ) );
  FDN1QM1P \Queue_reg[2][28]  ( .D(n502), .CPN(Clk_r), .Q(\Queue[2][28] ) );
  FDN1QM1P \Queue_reg[4][27]  ( .D(n405), .CPN(Clk_r), .Q(\Queue[4][27] ) );
  FDN1QM1P \Queue_reg[3][27]  ( .D(n533), .CPN(Clk_r), .Q(\Queue[3][27] ) );
  FDN1QM1P \Queue_reg[2][27]  ( .D(n501), .CPN(Clk_r), .Q(\Queue[2][27] ) );
  FDN1QM1P \Queue_reg[4][26]  ( .D(n404), .CPN(Clk_r), .Q(\Queue[4][26] ) );
  FDN1QM1P \Queue_reg[3][26]  ( .D(n532), .CPN(Clk_r), .Q(\Queue[3][26] ) );
  FDN1QM1P \Queue_reg[2][26]  ( .D(n500), .CPN(Clk_r), .Q(\Queue[2][26] ) );
  FDN1QM1P \Queue_reg[4][25]  ( .D(n403), .CPN(Clk_r), .Q(\Queue[4][25] ) );
  FDN1QM1P \Queue_reg[3][25]  ( .D(n531), .CPN(Clk_r), .Q(\Queue[3][25] ) );
  FDN1QM1P \Queue_reg[2][25]  ( .D(n499), .CPN(Clk_r), .Q(\Queue[2][25] ) );
  FDN1QM1P \Queue_reg[4][24]  ( .D(n402), .CPN(Clk_r), .Q(\Queue[4][24] ) );
  FDN1QM1P \Queue_reg[3][24]  ( .D(n530), .CPN(Clk_r), .Q(\Queue[3][24] ) );
  FDN1QM1P \Queue_reg[2][24]  ( .D(n498), .CPN(Clk_r), .Q(\Queue[2][24] ) );
  FDN1QM1P \Queue_reg[4][23]  ( .D(n401), .CPN(Clk_r), .Q(\Queue[4][23] ) );
  FDN1QM1P \Queue_reg[3][23]  ( .D(n529), .CPN(Clk_r), .Q(\Queue[3][23] ) );
  FDN1QM1P \Queue_reg[2][23]  ( .D(n497), .CPN(Clk_r), .Q(\Queue[2][23] ) );
  FDN1QM1P \Queue_reg[4][22]  ( .D(n400), .CPN(Clk_r), .Q(\Queue[4][22] ) );
  FDN1QM1P \Queue_reg[3][22]  ( .D(n528), .CPN(Clk_r), .Q(\Queue[3][22] ) );
  FDN1QM1P \Queue_reg[2][22]  ( .D(n496), .CPN(Clk_r), .Q(\Queue[2][22] ) );
  FDN1QM1P \Queue_reg[4][21]  ( .D(n399), .CPN(Clk_r), .Q(\Queue[4][21] ) );
  FDN1QM1P \Queue_reg[3][21]  ( .D(n527), .CPN(Clk_r), .Q(\Queue[3][21] ) );
  FDN1QM1P \Queue_reg[2][21]  ( .D(n495), .CPN(Clk_r), .Q(\Queue[2][21] ) );
  FDN1QM1P \Queue_reg[4][20]  ( .D(n398), .CPN(Clk_r), .Q(\Queue[4][20] ) );
  FDN1QM1P \Queue_reg[3][20]  ( .D(n526), .CPN(Clk_r), .Q(\Queue[3][20] ) );
  FDN1QM1P \Queue_reg[2][20]  ( .D(n494), .CPN(Clk_r), .Q(\Queue[2][20] ) );
  FDN1QM1P \Queue_reg[4][19]  ( .D(n397), .CPN(Clk_r), .Q(\Queue[4][19] ) );
  FDN1QM1P \Queue_reg[3][19]  ( .D(n525), .CPN(Clk_r), .Q(\Queue[3][19] ) );
  FDN1QM1P \Queue_reg[2][19]  ( .D(n493), .CPN(Clk_r), .Q(\Queue[2][19] ) );
  FDN1QM1P \Queue_reg[4][18]  ( .D(n396), .CPN(Clk_r), .Q(\Queue[4][18] ) );
  FDN1QM1P \Queue_reg[3][18]  ( .D(n524), .CPN(Clk_r), .Q(\Queue[3][18] ) );
  FDN1QM1P \Queue_reg[2][18]  ( .D(n492), .CPN(Clk_r), .Q(\Queue[2][18] ) );
  FDN1QM1P \Queue_reg[4][17]  ( .D(n395), .CPN(Clk_r), .Q(\Queue[4][17] ) );
  FDN1QM1P \Queue_reg[3][17]  ( .D(n523), .CPN(Clk_r), .Q(\Queue[3][17] ) );
  FDN1QM1P \Queue_reg[2][17]  ( .D(n491), .CPN(Clk_r), .Q(\Queue[2][17] ) );
  FDN1QM1P \Queue_reg[4][16]  ( .D(n394), .CPN(Clk_r), .Q(\Queue[4][16] ) );
  FDN1QM1P \Queue_reg[3][16]  ( .D(n522), .CPN(Clk_r), .Q(\Queue[3][16] ) );
  FDN1QM1P \Queue_reg[2][16]  ( .D(n490), .CPN(Clk_r), .Q(\Queue[2][16] ) );
  FDN1QM1P \Queue_reg[4][15]  ( .D(n393), .CPN(Clk_r), .Q(\Queue[4][15] ) );
  FDN1QM1P \Queue_reg[3][15]  ( .D(n521), .CPN(Clk_r), .Q(\Queue[3][15] ) );
  FDN1QM1P \Queue_reg[2][15]  ( .D(n489), .CPN(Clk_r), .Q(\Queue[2][15] ) );
  FDN1QM1P \Queue_reg[4][14]  ( .D(n392), .CPN(Clk_r), .Q(\Queue[4][14] ) );
  FDN1QM1P \Queue_reg[3][14]  ( .D(n520), .CPN(Clk_r), .Q(\Queue[3][14] ) );
  FDN1QM1P \Queue_reg[2][14]  ( .D(n488), .CPN(Clk_r), .Q(\Queue[2][14] ) );
  FDN1QM1P \Queue_reg[4][13]  ( .D(n391), .CPN(Clk_r), .Q(\Queue[4][13] ) );
  FDN1QM1P \Queue_reg[3][13]  ( .D(n519), .CPN(Clk_r), .Q(\Queue[3][13] ) );
  FDN1QM1P \Queue_reg[2][13]  ( .D(n487), .CPN(Clk_r), .Q(\Queue[2][13] ) );
  FDN1QM1P \Queue_reg[4][12]  ( .D(n390), .CPN(Clk_r), .Q(\Queue[4][12] ) );
  FDN1QM1P \Queue_reg[3][12]  ( .D(n518), .CPN(Clk_r), .Q(\Queue[3][12] ) );
  FDN1QM1P \Queue_reg[2][12]  ( .D(n486), .CPN(Clk_r), .Q(\Queue[2][12] ) );
  FDN1QM1P \Queue_reg[4][11]  ( .D(n389), .CPN(Clk_r), .Q(\Queue[4][11] ) );
  FDN1QM1P \Queue_reg[3][11]  ( .D(n517), .CPN(Clk_r), .Q(\Queue[3][11] ) );
  FDN1QM1P \Queue_reg[2][11]  ( .D(n485), .CPN(Clk_r), .Q(\Queue[2][11] ) );
  FDN1QM1P \Queue_reg[4][10]  ( .D(n388), .CPN(Clk_r), .Q(\Queue[4][10] ) );
  FDN1QM1P \Queue_reg[3][10]  ( .D(n516), .CPN(Clk_r), .Q(\Queue[3][10] ) );
  FDN1QM1P \Queue_reg[2][10]  ( .D(n484), .CPN(Clk_r), .Q(\Queue[2][10] ) );
  FDN1QM1P \Queue_reg[4][9]  ( .D(n387), .CPN(Clk_r), .Q(\Queue[4][9] ) );
  FDN1QM1P \Queue_reg[3][9]  ( .D(n515), .CPN(Clk_r), .Q(\Queue[3][9] ) );
  FDN1QM1P \Queue_reg[2][9]  ( .D(n483), .CPN(Clk_r), .Q(\Queue[2][9] ) );
  FDN1QM1P \Queue_reg[4][8]  ( .D(n386), .CPN(Clk_r), .Q(\Queue[4][8] ) );
  FDN1QM1P \Queue_reg[3][8]  ( .D(n514), .CPN(Clk_r), .Q(\Queue[3][8] ) );
  FDN1QM1P \Queue_reg[2][8]  ( .D(n482), .CPN(Clk_r), .Q(\Queue[2][8] ) );
  FDN1QM1P \Queue_reg[4][7]  ( .D(n385), .CPN(Clk_r), .Q(\Queue[4][7] ) );
  FDN1QM1P \Queue_reg[3][7]  ( .D(n513), .CPN(Clk_r), .Q(\Queue[3][7] ) );
  FDN1QM1P \Queue_reg[2][7]  ( .D(n481), .CPN(Clk_r), .Q(\Queue[2][7] ) );
  FDN1QM1P \Queue_reg[4][6]  ( .D(n384), .CPN(Clk_r), .Q(\Queue[4][6] ) );
  FDN1QM1P \Queue_reg[3][6]  ( .D(n512), .CPN(Clk_r), .Q(\Queue[3][6] ) );
  FDN1QM1P \Queue_reg[2][6]  ( .D(n480), .CPN(Clk_r), .Q(\Queue[2][6] ) );
  FDN1QM1P \Queue_reg[4][5]  ( .D(n383), .CPN(Clk_r), .Q(\Queue[4][5] ) );
  FDN1QM1P \Queue_reg[3][5]  ( .D(n511), .CPN(Clk_r), .Q(\Queue[3][5] ) );
  FDN1QM1P \Queue_reg[2][5]  ( .D(n479), .CPN(Clk_r), .Q(\Queue[2][5] ) );
  FDN1QM1P \Queue_reg[4][4]  ( .D(n382), .CPN(Clk_r), .Q(\Queue[4][4] ) );
  FDN1QM1P \Queue_reg[3][4]  ( .D(n510), .CPN(Clk_r), .Q(\Queue[3][4] ) );
  FDN1QM1P \Queue_reg[2][4]  ( .D(n478), .CPN(Clk_r), .Q(\Queue[2][4] ) );
  FDN1QM1P \Queue_reg[4][3]  ( .D(n381), .CPN(Clk_r), .Q(\Queue[4][3] ) );
  FDN1QM1P \Queue_reg[3][3]  ( .D(n509), .CPN(Clk_r), .Q(\Queue[3][3] ) );
  FDN1QM1P \Queue_reg[2][3]  ( .D(n477), .CPN(Clk_r), .Q(\Queue[2][3] ) );
  FDN1QM1P \Queue_reg[4][2]  ( .D(n380), .CPN(Clk_r), .Q(\Queue[4][2] ) );
  FDN1QM1P \Queue_reg[3][2]  ( .D(n508), .CPN(Clk_r), .Q(\Queue[3][2] ) );
  FDN1QM1P \Queue_reg[2][2]  ( .D(n476), .CPN(Clk_r), .Q(\Queue[2][2] ) );
  FDN1QM1P \Queue_reg[4][1]  ( .D(n379), .CPN(Clk_r), .Q(\Queue[4][1] ) );
  FDN1QM1P \Queue_reg[3][1]  ( .D(n507), .CPN(Clk_r), .Q(\Queue[3][1] ) );
  FDN1QM1P \Queue_reg[2][1]  ( .D(n475), .CPN(Clk_r), .Q(\Queue[2][1] ) );
  FDN1QM1P \Queue_reg[4][0]  ( .D(n378), .CPN(Clk_r), .Q(\Queue[4][0] ) );
  FDN1QM1P \Queue_reg[3][0]  ( .D(n506), .CPN(Clk_r), .Q(\Queue[3][0] ) );
  FDN1QM1P \Queue_reg[2][0]  ( .D(n474), .CPN(Clk_r), .Q(\Queue[2][0] ) );
  FDN1QM1P \Queue_reg[4][31]  ( .D(n377), .CPN(Clk_r), .Q(\Queue[4][31] ) );
  FDN1QM1P \Queue_reg[3][31]  ( .D(n537), .CPN(Clk_r), .Q(\Queue[3][31] ) );
  FDN1QM1P \Queue_reg[2][31]  ( .D(n505), .CPN(Clk_r), .Q(\Queue[2][31] ) );
  FDN2QM1P Full_reg ( .D(n409), .CPN(Clk_r), .CD(Rst_n), .Q(Full) );
  FDN1QM1P \Queue_reg[1][31]  ( .D(n441), .CPN(Clk_r), .Q(\Queue[1][31] ) );
  FDN1QM1P \Queue_reg[0][31]  ( .D(n473), .CPN(Clk_r), .Q(Packet_Out[31]) );
  FDN1QM1P \Queue_reg[1][30]  ( .D(n440), .CPN(Clk_r), .Q(\Queue[1][30] ) );
  FDN1QM1P \Queue_reg[0][30]  ( .D(n472), .CPN(Clk_r), .Q(Packet_Out[30]) );
  FDN1QM1P \Queue_reg[1][29]  ( .D(n439), .CPN(Clk_r), .Q(\Queue[1][29] ) );
  FDN1QM1P \Queue_reg[0][29]  ( .D(n471), .CPN(Clk_r), .Q(Packet_Out[29]) );
  FDN1QM1P \Queue_reg[1][28]  ( .D(n438), .CPN(Clk_r), .Q(\Queue[1][28] ) );
  FDN1QM1P \Queue_reg[0][28]  ( .D(n470), .CPN(Clk_r), .Q(Packet_Out[28]) );
  FDN1QM1P \Queue_reg[1][27]  ( .D(n437), .CPN(Clk_r), .Q(\Queue[1][27] ) );
  FDN1QM1P \Queue_reg[0][27]  ( .D(n469), .CPN(Clk_r), .Q(Packet_Out[27]) );
  FDN1QM1P \Queue_reg[1][26]  ( .D(n436), .CPN(Clk_r), .Q(\Queue[1][26] ) );
  FDN1QM1P \Queue_reg[0][26]  ( .D(n468), .CPN(Clk_r), .Q(Packet_Out[26]) );
  FDN1QM1P \Queue_reg[1][25]  ( .D(n435), .CPN(Clk_r), .Q(\Queue[1][25] ) );
  FDN1QM1P \Queue_reg[0][25]  ( .D(n467), .CPN(Clk_r), .Q(Packet_Out[25]) );
  FDN1QM1P \Queue_reg[1][24]  ( .D(n434), .CPN(Clk_r), .Q(\Queue[1][24] ) );
  FDN1QM1P \Queue_reg[0][24]  ( .D(n466), .CPN(Clk_r), .Q(Packet_Out[24]) );
  FDN1QM1P \Queue_reg[1][23]  ( .D(n433), .CPN(Clk_r), .Q(\Queue[1][23] ) );
  FDN1QM1P \Queue_reg[0][23]  ( .D(n465), .CPN(Clk_r), .Q(Packet_Out[23]) );
  FDN1QM1P \Queue_reg[1][22]  ( .D(n432), .CPN(Clk_r), .Q(\Queue[1][22] ) );
  FDN1QM1P \Queue_reg[0][22]  ( .D(n464), .CPN(Clk_r), .Q(Packet_Out[22]) );
  FDN1QM1P \Queue_reg[1][21]  ( .D(n431), .CPN(Clk_r), .Q(\Queue[1][21] ) );
  FDN1QM1P \Queue_reg[0][21]  ( .D(n463), .CPN(Clk_r), .Q(Packet_Out[21]) );
  FDN1QM1P \Queue_reg[1][20]  ( .D(n430), .CPN(Clk_r), .Q(\Queue[1][20] ) );
  FDN1QM1P \Queue_reg[0][20]  ( .D(n462), .CPN(Clk_r), .Q(Packet_Out[20]) );
  FDN1QM1P \Queue_reg[1][19]  ( .D(n429), .CPN(Clk_r), .Q(\Queue[1][19] ) );
  FDN1QM1P \Queue_reg[0][19]  ( .D(n461), .CPN(Clk_r), .Q(Packet_Out[19]) );
  FDN1QM1P \Queue_reg[1][18]  ( .D(n428), .CPN(Clk_r), .Q(\Queue[1][18] ) );
  FDN1QM1P \Queue_reg[0][18]  ( .D(n460), .CPN(Clk_r), .Q(Packet_Out[18]) );
  FDN1QM1P \Queue_reg[1][17]  ( .D(n427), .CPN(Clk_r), .Q(\Queue[1][17] ) );
  FDN1QM1P \Queue_reg[0][17]  ( .D(n459), .CPN(Clk_r), .Q(Packet_Out[17]) );
  FDN1QM1P \Queue_reg[1][16]  ( .D(n426), .CPN(Clk_r), .Q(\Queue[1][16] ) );
  FDN1QM1P \Queue_reg[0][16]  ( .D(n458), .CPN(Clk_r), .Q(Packet_Out[16]) );
  FDN1QM1P \Queue_reg[1][15]  ( .D(n425), .CPN(Clk_r), .Q(\Queue[1][15] ) );
  FDN1QM1P \Queue_reg[0][15]  ( .D(n457), .CPN(Clk_r), .Q(Packet_Out[15]) );
  FDN1QM1P \Queue_reg[1][14]  ( .D(n424), .CPN(Clk_r), .Q(\Queue[1][14] ) );
  FDN1QM1P \Queue_reg[0][14]  ( .D(n456), .CPN(Clk_r), .Q(Packet_Out[14]) );
  FDN1QM1P \Queue_reg[1][13]  ( .D(n423), .CPN(Clk_r), .Q(\Queue[1][13] ) );
  FDN1QM1P \Queue_reg[0][13]  ( .D(n455), .CPN(Clk_r), .Q(Packet_Out[13]) );
  FDN1QM1P \Queue_reg[1][12]  ( .D(n422), .CPN(Clk_r), .Q(\Queue[1][12] ) );
  FDN1QM1P \Queue_reg[0][12]  ( .D(n454), .CPN(Clk_r), .Q(Packet_Out[12]) );
  FDN1QM1P \Queue_reg[1][11]  ( .D(n421), .CPN(Clk_r), .Q(\Queue[1][11] ) );
  FDN1QM1P \Queue_reg[0][11]  ( .D(n453), .CPN(Clk_r), .Q(Packet_Out[11]) );
  FDN1QM1P \Queue_reg[1][10]  ( .D(n420), .CPN(Clk_r), .Q(\Queue[1][10] ) );
  FDN1QM1P \Queue_reg[0][10]  ( .D(n452), .CPN(Clk_r), .Q(Packet_Out[10]) );
  FDN1QM1P \Queue_reg[1][9]  ( .D(n419), .CPN(Clk_r), .Q(\Queue[1][9] ) );
  FDN1QM1P \Queue_reg[0][9]  ( .D(n451), .CPN(Clk_r), .Q(Packet_Out[9]) );
  FDN1QM1P \Queue_reg[1][8]  ( .D(n418), .CPN(Clk_r), .Q(\Queue[1][8] ) );
  FDN1QM1P \Queue_reg[0][8]  ( .D(n450), .CPN(Clk_r), .Q(Packet_Out[8]) );
  FDN1QM1P \Queue_reg[1][7]  ( .D(n417), .CPN(Clk_r), .Q(\Queue[1][7] ) );
  FDN1QM1P \Queue_reg[0][7]  ( .D(n449), .CPN(Clk_r), .Q(Packet_Out[7]) );
  FDN1QM1P \Queue_reg[1][6]  ( .D(n416), .CPN(Clk_r), .Q(\Queue[1][6] ) );
  FDN1QM1P \Queue_reg[0][6]  ( .D(n448), .CPN(Clk_r), .Q(Packet_Out[6]) );
  FDN1QM1P \Queue_reg[1][5]  ( .D(n415), .CPN(Clk_r), .Q(\Queue[1][5] ) );
  FDN1QM1P \Queue_reg[0][5]  ( .D(n447), .CPN(Clk_r), .Q(Packet_Out[5]) );
  FDN1QM1P \Queue_reg[1][4]  ( .D(n414), .CPN(Clk_r), .Q(\Queue[1][4] ) );
  FDN1QM1P \Queue_reg[0][4]  ( .D(n446), .CPN(Clk_r), .Q(Packet_Out[4]) );
  FDN1QM1P \Queue_reg[1][3]  ( .D(n413), .CPN(Clk_r), .Q(\Queue[1][3] ) );
  FDN1QM1P \Queue_reg[0][3]  ( .D(n445), .CPN(Clk_r), .Q(Packet_Out[3]) );
  FDN1QM1P \Queue_reg[1][2]  ( .D(n412), .CPN(Clk_r), .Q(\Queue[1][2] ) );
  FDN1QM1P \Queue_reg[0][2]  ( .D(n444), .CPN(Clk_r), .Q(Packet_Out[2]) );
  FDN1QM1P \Queue_reg[1][1]  ( .D(n411), .CPN(Clk_r), .Q(\Queue[1][1] ) );
  FDN1QM1P \Queue_reg[0][1]  ( .D(n443), .CPN(Clk_r), .Q(Packet_Out[1]) );
  FDN1QM1P \Queue_reg[1][0]  ( .D(n410), .CPN(Clk_r), .Q(\Queue[1][0] ) );
  FDN1QM1P \Queue_reg[0][0]  ( .D(n442), .CPN(Clk_r), .Q(Packet_Out[0]) );
  FDN2QM1P Empty_reg ( .D(n539), .CPN(Clk_r), .CD(Rst_n), .Q(n538) );
  BUFM1P U3 ( .A(n130), .Z(n7) );
  BUFM1P U4 ( .A(n203), .Z(n9) );
  BUFM2P U5 ( .A(n130), .Z(n6) );
  BUFM2P U6 ( .A(n203), .Z(n8) );
  NR2FM1P U7 ( .A(Read_Ack), .B(n96), .Z(n15) );
  N1M1P U8 ( .A(Read_Ack), .Z(n134) );
  BUFM3P U9 ( .A(n53), .Z(n3) );
  OAI211M4P U10 ( .A(n97), .B(n134), .C(Write_Ack), .D(n21), .Z(n56) );
  OAI211M4P U11 ( .A(n137), .B(n134), .C(Write_Ack), .D(n95), .Z(n132) );
  OAI211M4P U12 ( .A(n139), .B(n134), .C(Write_Ack), .D(n133), .Z(n205) );
  AOI21M3P U13 ( .A(Write_Ack), .B(n139), .C(n138), .Z(n202) );
  AOI21M3P U14 ( .A(Write_Ack), .B(n137), .C(n138), .Z(n129) );
  N1M2P U15 ( .A(n59), .Z(n91) );
  OAI211M4P U16 ( .A(n373), .B(n134), .C(Write_Ack), .D(n59), .Z(n94) );
  NR2FM3P U17 ( .A(n58), .B(n18), .Z(n17) );
  N1M1P U18 ( .A(n139), .Z(n18) );
  NR3M1P U19 ( .A(Count[0]), .B(Count[1]), .C(n16), .Z(n139) );
  NR3M1P U20 ( .A(n20), .B(Count[2]), .C(Count[1]), .Z(n373) );
  NR3M1P U21 ( .A(Count[0]), .B(Count[2]), .C(n19), .Z(n97) );
  NR3M1P U22 ( .A(Count[2]), .B(n20), .C(n19), .Z(n137) );
  N1M1P U23 ( .A(Count[1]), .Z(n19) );
  N1M1P U24 ( .A(Count[2]), .Z(n16) );
  N1M1P U25 ( .A(Count[0]), .Z(n20) );
  ND2M2P U26 ( .A(n15), .B(Rst_n), .Z(n58) );
  AOI21M6P U27 ( .A(Write_Ack), .B(n97), .C(n138), .Z(n54) );
  AOI21M6P U28 ( .A(Write_Ack), .B(n373), .C(n138), .Z(n92) );
  ND2M2P U29 ( .A(Read_Ack), .B(Rst_n), .Z(n138) );
  BUFM2P U30 ( .A(n91), .Z(n5) );
  BUFM2P U31 ( .A(n53), .Z(n4) );
  N1M2P U32 ( .A(n15), .Z(n136) );
  AOI22M1P U33 ( .A(\Queue[2][1] ), .B(n6), .C(n129), .D(\Queue[3][1] ), .Z(
        n99) );
  N1M1P U34 ( .A(n538), .Z(Empty) );
  OAI21M1P U35 ( .A(Write_Ack), .B(Read_Ack), .C(n21), .Z(n53) );
  N1M2P U36 ( .A(Write_Ack), .Z(n96) );
  OAI211M1P U37 ( .A(n137), .B(n136), .C(Rst_n), .D(n135), .Z(n203) );
  OAI211M1P U38 ( .A(n97), .B(n136), .C(Rst_n), .D(n135), .Z(n130) );
  NR2M1P U39 ( .A(n134), .B(Write_Ack), .Z(n208) );
  NR2M1P U40 ( .A(n15), .B(n208), .Z(n207) );
  AOI22CDNM1P U41 ( .A(n207), .B(n20), .C(n207), .D(n20), .Z(n374) );
  N1M1P U42 ( .A(n208), .Z(n14) );
  AOI22M1P U43 ( .A(Count[0]), .B(n136), .C(n14), .D(n20), .Z(n11) );
  AOI22CDNM1P U44 ( .A(Count[1]), .B(n11), .C(n11), .D(Count[1]), .Z(n375) );
  ND3M1P U45 ( .A(n20), .B(n16), .C(n19), .Z(n57) );
  ND2M1P U46 ( .A(Count[1]), .B(Read_Ack), .Z(n10) );
  OAI211M1P U47 ( .A(Count[1]), .B(n136), .C(n11), .D(n10), .Z(n12) );
  AOI22M1P U48 ( .A(n15), .B(n137), .C(Count[2]), .D(n12), .Z(n13) );
  OAI21M1P U49 ( .A(n57), .B(n14), .C(n13), .Z(n376) );
  N1M1P U50 ( .A(Packet_In[31]), .Z(n206) );
  AOI22CDNM1P U51 ( .A(n17), .B(n206), .C(\Queue[4][31] ), .D(n17), .Z(n377)
         );
  N1M1P U52 ( .A(Packet_In[0]), .Z(n141) );
  AOI22CDNM1P U53 ( .A(n17), .B(n141), .C(\Queue[4][0] ), .D(n17), .Z(n378) );
  N1M1P U54 ( .A(Packet_In[1]), .Z(n143) );
  AOI22CDNM1P U55 ( .A(n17), .B(n143), .C(\Queue[4][1] ), .D(n17), .Z(n379) );
  N1M1P U56 ( .A(Packet_In[2]), .Z(n145) );
  AOI22CDNM1P U57 ( .A(n17), .B(n145), .C(\Queue[4][2] ), .D(n17), .Z(n380) );
  N1M1P U58 ( .A(Packet_In[3]), .Z(n147) );
  AOI22CDNM1P U59 ( .A(n17), .B(n147), .C(\Queue[4][3] ), .D(n17), .Z(n381) );
  N1M1P U60 ( .A(Packet_In[4]), .Z(n149) );
  AOI22CDNM1P U61 ( .A(n17), .B(n149), .C(\Queue[4][4] ), .D(n17), .Z(n382) );
  N1M1P U62 ( .A(Packet_In[5]), .Z(n151) );
  AOI22CDNM1P U63 ( .A(n17), .B(n151), .C(\Queue[4][5] ), .D(n17), .Z(n383) );
  N1M1P U64 ( .A(Packet_In[6]), .Z(n153) );
  AOI22CDNM1P U65 ( .A(n17), .B(n153), .C(\Queue[4][6] ), .D(n17), .Z(n384) );
  N1M1P U66 ( .A(Packet_In[7]), .Z(n155) );
  AOI22CDNM1P U67 ( .A(n17), .B(n155), .C(\Queue[4][7] ), .D(n17), .Z(n385) );
  N1M1P U68 ( .A(Packet_In[8]), .Z(n157) );
  AOI22CDNM1P U69 ( .A(n17), .B(n157), .C(\Queue[4][8] ), .D(n17), .Z(n386) );
  N1M1P U70 ( .A(Packet_In[9]), .Z(n159) );
  AOI22CDNM1P U71 ( .A(n17), .B(n159), .C(\Queue[4][9] ), .D(n17), .Z(n387) );
  N1M1P U72 ( .A(Packet_In[10]), .Z(n161) );
  AOI22CDNM1P U73 ( .A(n17), .B(n161), .C(\Queue[4][10] ), .D(n17), .Z(n388)
         );
  N1M1P U74 ( .A(Packet_In[11]), .Z(n163) );
  AOI22CDNM1P U75 ( .A(n17), .B(n163), .C(\Queue[4][11] ), .D(n17), .Z(n389)
         );
  N1M1P U76 ( .A(Packet_In[12]), .Z(n165) );
  AOI22CDNM1P U77 ( .A(n17), .B(n165), .C(\Queue[4][12] ), .D(n17), .Z(n390)
         );
  N1M1P U78 ( .A(Packet_In[13]), .Z(n167) );
  AOI22CDNM1P U79 ( .A(n17), .B(n167), .C(\Queue[4][13] ), .D(n17), .Z(n391)
         );
  N1M1P U80 ( .A(Packet_In[14]), .Z(n169) );
  AOI22CDNM1P U81 ( .A(n17), .B(n169), .C(\Queue[4][14] ), .D(n17), .Z(n392)
         );
  N1M1P U82 ( .A(Packet_In[15]), .Z(n171) );
  AOI22CDNM1P U83 ( .A(n17), .B(n171), .C(\Queue[4][15] ), .D(n17), .Z(n393)
         );
  N1M1P U84 ( .A(Packet_In[16]), .Z(n173) );
  AOI22CDNM1P U85 ( .A(n17), .B(n173), .C(\Queue[4][16] ), .D(n17), .Z(n394)
         );
  N1M1P U86 ( .A(Packet_In[17]), .Z(n175) );
  AOI22CDNM1P U87 ( .A(n17), .B(n175), .C(\Queue[4][17] ), .D(n17), .Z(n395)
         );
  N1M1P U88 ( .A(Packet_In[18]), .Z(n177) );
  AOI22CDNM1P U89 ( .A(n17), .B(n177), .C(\Queue[4][18] ), .D(n17), .Z(n396)
         );
  N1M1P U90 ( .A(Packet_In[19]), .Z(n179) );
  AOI22CDNM1P U91 ( .A(n17), .B(n179), .C(\Queue[4][19] ), .D(n17), .Z(n397)
         );
  N1M1P U92 ( .A(Packet_In[20]), .Z(n181) );
  AOI22CDNM1P U93 ( .A(n17), .B(n181), .C(\Queue[4][20] ), .D(n17), .Z(n398)
         );
  N1M1P U94 ( .A(Packet_In[21]), .Z(n183) );
  AOI22CDNM1P U95 ( .A(n17), .B(n183), .C(\Queue[4][21] ), .D(n17), .Z(n399)
         );
  N1M1P U96 ( .A(Packet_In[22]), .Z(n185) );
  AOI22CDNM1P U97 ( .A(n17), .B(n185), .C(\Queue[4][22] ), .D(n17), .Z(n400)
         );
  N1M1P U98 ( .A(Packet_In[23]), .Z(n187) );
  AOI22CDNM1P U99 ( .A(n17), .B(n187), .C(\Queue[4][23] ), .D(n17), .Z(n401)
         );
  N1M1P U100 ( .A(Packet_In[24]), .Z(n189) );
  AOI22CDNM1P U101 ( .A(n17), .B(n189), .C(\Queue[4][24] ), .D(n17), .Z(n402)
         );
  N1M1P U102 ( .A(Packet_In[25]), .Z(n191) );
  AOI22CDNM1P U103 ( .A(n17), .B(n191), .C(\Queue[4][25] ), .D(n17), .Z(n403)
         );
  N1M1P U104 ( .A(Packet_In[26]), .Z(n193) );
  AOI22CDNM1P U105 ( .A(n17), .B(n193), .C(\Queue[4][26] ), .D(n17), .Z(n404)
         );
  N1M1P U106 ( .A(Packet_In[27]), .Z(n195) );
  AOI22CDNM1P U107 ( .A(n17), .B(n195), .C(\Queue[4][27] ), .D(n17), .Z(n405)
         );
  N1M1P U108 ( .A(Packet_In[28]), .Z(n197) );
  AOI22CDNM1P U109 ( .A(n17), .B(n197), .C(\Queue[4][28] ), .D(n17), .Z(n406)
         );
  N1M1P U110 ( .A(Packet_In[29]), .Z(n199) );
  AOI22CDNM1P U111 ( .A(n17), .B(n199), .C(\Queue[4][29] ), .D(n17), .Z(n407)
         );
  N1M1P U112 ( .A(Packet_In[30]), .Z(n201) );
  AOI22CDNM1P U113 ( .A(n17), .B(n201), .C(\Queue[4][30] ), .D(n17), .Z(n408)
         );
  OAI22CDNM1P U114 ( .A(n136), .B(n18), .C(n207), .D(Full), .Z(n409) );
  OA21M1P U115 ( .A(n136), .B(n373), .C(Rst_n), .Z(n21) );
  AOI22M1P U116 ( .A(\Queue[2][0] ), .B(n54), .C(\Queue[1][0] ), .D(n53), .Z(
        n22) );
  OAI21M1P U117 ( .A(n141), .B(n56), .C(n22), .Z(n410) );
  AOI22M1P U118 ( .A(n54), .B(\Queue[2][1] ), .C(\Queue[1][1] ), .D(n53), .Z(
        n23) );
  OAI21M1P U119 ( .A(n56), .B(n143), .C(n23), .Z(n411) );
  AOI22M1P U120 ( .A(n54), .B(\Queue[2][2] ), .C(\Queue[1][2] ), .D(n53), .Z(
        n24) );
  OAI21M1P U121 ( .A(n56), .B(n145), .C(n24), .Z(n412) );
  AOI22M1P U122 ( .A(n54), .B(\Queue[2][3] ), .C(\Queue[1][3] ), .D(n3), .Z(
        n25) );
  OAI21M1P U123 ( .A(n56), .B(n147), .C(n25), .Z(n413) );
  AOI22M1P U124 ( .A(n54), .B(\Queue[2][4] ), .C(\Queue[1][4] ), .D(n4), .Z(
        n26) );
  OAI21M1P U125 ( .A(n56), .B(n149), .C(n26), .Z(n414) );
  AOI22M1P U126 ( .A(n54), .B(\Queue[2][5] ), .C(\Queue[1][5] ), .D(n3), .Z(
        n27) );
  OAI21M1P U127 ( .A(n56), .B(n151), .C(n27), .Z(n415) );
  AOI22M1P U128 ( .A(n54), .B(\Queue[2][6] ), .C(\Queue[1][6] ), .D(n4), .Z(
        n28) );
  OAI21M1P U129 ( .A(n56), .B(n153), .C(n28), .Z(n416) );
  AOI22M1P U130 ( .A(n54), .B(\Queue[2][7] ), .C(\Queue[1][7] ), .D(n4), .Z(
        n29) );
  OAI21M1P U131 ( .A(n56), .B(n155), .C(n29), .Z(n417) );
  AOI22M1P U132 ( .A(n54), .B(\Queue[2][8] ), .C(\Queue[1][8] ), .D(n4), .Z(
        n30) );
  OAI21M1P U133 ( .A(n56), .B(n157), .C(n30), .Z(n418) );
  AOI22M1P U134 ( .A(n54), .B(\Queue[2][9] ), .C(\Queue[1][9] ), .D(n3), .Z(
        n31) );
  OAI21M1P U135 ( .A(n56), .B(n159), .C(n31), .Z(n419) );
  AOI22M1P U136 ( .A(n54), .B(\Queue[2][10] ), .C(\Queue[1][10] ), .D(n3), .Z(
        n32) );
  OAI21M1P U137 ( .A(n56), .B(n161), .C(n32), .Z(n420) );
  AOI22M1P U138 ( .A(n54), .B(\Queue[2][11] ), .C(\Queue[1][11] ), .D(n3), .Z(
        n33) );
  OAI21M1P U139 ( .A(n56), .B(n163), .C(n33), .Z(n421) );
  AOI22M1P U140 ( .A(n54), .B(\Queue[2][12] ), .C(\Queue[1][12] ), .D(n3), .Z(
        n34) );
  OAI21M1P U141 ( .A(n56), .B(n165), .C(n34), .Z(n422) );
  AOI22M1P U142 ( .A(n54), .B(\Queue[2][13] ), .C(\Queue[1][13] ), .D(n3), .Z(
        n35) );
  OAI21M1P U143 ( .A(n56), .B(n167), .C(n35), .Z(n423) );
  AOI22M1P U144 ( .A(n54), .B(\Queue[2][14] ), .C(\Queue[1][14] ), .D(n3), .Z(
        n36) );
  OAI21M1P U145 ( .A(n56), .B(n169), .C(n36), .Z(n424) );
  AOI22M1P U146 ( .A(n54), .B(\Queue[2][15] ), .C(\Queue[1][15] ), .D(n3), .Z(
        n37) );
  OAI21M1P U147 ( .A(n56), .B(n171), .C(n37), .Z(n425) );
  AOI22M1P U148 ( .A(n54), .B(\Queue[2][16] ), .C(\Queue[1][16] ), .D(n3), .Z(
        n38) );
  OAI21M1P U149 ( .A(n56), .B(n173), .C(n38), .Z(n426) );
  AOI22M1P U150 ( .A(n54), .B(\Queue[2][17] ), .C(\Queue[1][17] ), .D(n3), .Z(
        n39) );
  OAI21M1P U151 ( .A(n56), .B(n175), .C(n39), .Z(n427) );
  AOI22M1P U152 ( .A(n54), .B(\Queue[2][18] ), .C(\Queue[1][18] ), .D(n4), .Z(
        n40) );
  OAI21M1P U153 ( .A(n56), .B(n177), .C(n40), .Z(n428) );
  AOI22M1P U154 ( .A(n54), .B(\Queue[2][19] ), .C(\Queue[1][19] ), .D(n4), .Z(
        n41) );
  OAI21M1P U155 ( .A(n56), .B(n179), .C(n41), .Z(n429) );
  AOI22M1P U156 ( .A(n54), .B(\Queue[2][20] ), .C(\Queue[1][20] ), .D(n4), .Z(
        n42) );
  OAI21M1P U157 ( .A(n56), .B(n181), .C(n42), .Z(n430) );
  AOI22M1P U158 ( .A(n54), .B(\Queue[2][21] ), .C(\Queue[1][21] ), .D(n4), .Z(
        n43) );
  OAI21M1P U159 ( .A(n56), .B(n183), .C(n43), .Z(n431) );
  AOI22M1P U160 ( .A(n54), .B(\Queue[2][22] ), .C(\Queue[1][22] ), .D(n4), .Z(
        n44) );
  OAI21M1P U161 ( .A(n56), .B(n185), .C(n44), .Z(n432) );
  AOI22M1P U162 ( .A(n54), .B(\Queue[2][23] ), .C(\Queue[1][23] ), .D(n4), .Z(
        n45) );
  OAI21M1P U163 ( .A(n56), .B(n187), .C(n45), .Z(n433) );
  AOI22M1P U164 ( .A(n54), .B(\Queue[2][24] ), .C(\Queue[1][24] ), .D(n4), .Z(
        n46) );
  OAI21M1P U165 ( .A(n56), .B(n189), .C(n46), .Z(n434) );
  AOI22M1P U166 ( .A(n54), .B(\Queue[2][25] ), .C(\Queue[1][25] ), .D(n4), .Z(
        n47) );
  OAI21M1P U167 ( .A(n56), .B(n191), .C(n47), .Z(n435) );
  AOI22M1P U168 ( .A(n54), .B(\Queue[2][26] ), .C(\Queue[1][26] ), .D(n4), .Z(
        n48) );
  OAI21M1P U169 ( .A(n56), .B(n193), .C(n48), .Z(n436) );
  AOI22M1P U170 ( .A(n54), .B(\Queue[2][27] ), .C(\Queue[1][27] ), .D(n3), .Z(
        n49) );
  OAI21M1P U171 ( .A(n56), .B(n195), .C(n49), .Z(n437) );
  AOI22M1P U172 ( .A(n54), .B(\Queue[2][28] ), .C(\Queue[1][28] ), .D(n3), .Z(
        n50) );
  OAI21M1P U173 ( .A(n56), .B(n197), .C(n50), .Z(n438) );
  AOI22M1P U174 ( .A(n54), .B(\Queue[2][29] ), .C(\Queue[1][29] ), .D(n3), .Z(
        n51) );
  OAI21M1P U175 ( .A(n56), .B(n199), .C(n51), .Z(n439) );
  AOI22M1P U176 ( .A(n54), .B(\Queue[2][30] ), .C(\Queue[1][30] ), .D(n3), .Z(
        n52) );
  OAI21M1P U177 ( .A(n56), .B(n201), .C(n52), .Z(n440) );
  AOI22M1P U178 ( .A(n54), .B(\Queue[2][31] ), .C(\Queue[1][31] ), .D(n3), .Z(
        n55) );
  OAI21M1P U179 ( .A(n56), .B(n206), .C(n55), .Z(n441) );
  OAI21M1P U180 ( .A(n58), .B(n57), .C(n138), .Z(n59) );
  AOI22M1P U181 ( .A(\Queue[1][0] ), .B(n92), .C(n5), .D(Packet_Out[0]), .Z(
        n60) );
  OAI21M1P U182 ( .A(n141), .B(n94), .C(n60), .Z(n442) );
  AOI22M1P U183 ( .A(\Queue[1][1] ), .B(n92), .C(n91), .D(Packet_Out[1]), .Z(
        n61) );
  OAI21M1P U184 ( .A(n143), .B(n94), .C(n61), .Z(n443) );
  AOI22M1P U185 ( .A(\Queue[1][2] ), .B(n92), .C(n91), .D(Packet_Out[2]), .Z(
        n62) );
  OAI21M1P U186 ( .A(n145), .B(n94), .C(n62), .Z(n444) );
  AOI22M1P U187 ( .A(\Queue[1][3] ), .B(n92), .C(n91), .D(Packet_Out[3]), .Z(
        n63) );
  OAI21M1P U188 ( .A(n147), .B(n94), .C(n63), .Z(n445) );
  AOI22M1P U189 ( .A(\Queue[1][4] ), .B(n92), .C(n91), .D(Packet_Out[4]), .Z(
        n64) );
  OAI21M1P U190 ( .A(n149), .B(n94), .C(n64), .Z(n446) );
  AOI22M1P U191 ( .A(\Queue[1][5] ), .B(n92), .C(n91), .D(Packet_Out[5]), .Z(
        n65) );
  OAI21M1P U192 ( .A(n151), .B(n94), .C(n65), .Z(n447) );
  AOI22M1P U193 ( .A(\Queue[1][6] ), .B(n92), .C(n91), .D(Packet_Out[6]), .Z(
        n66) );
  OAI21M1P U194 ( .A(n153), .B(n94), .C(n66), .Z(n448) );
  AOI22M1P U195 ( .A(\Queue[1][7] ), .B(n92), .C(n91), .D(Packet_Out[7]), .Z(
        n67) );
  OAI21M1P U196 ( .A(n155), .B(n94), .C(n67), .Z(n449) );
  AOI22M1P U197 ( .A(\Queue[1][8] ), .B(n92), .C(n91), .D(Packet_Out[8]), .Z(
        n68) );
  OAI21M1P U198 ( .A(n157), .B(n94), .C(n68), .Z(n450) );
  AOI22M1P U199 ( .A(\Queue[1][9] ), .B(n92), .C(n91), .D(Packet_Out[9]), .Z(
        n69) );
  OAI21M1P U200 ( .A(n159), .B(n94), .C(n69), .Z(n451) );
  AOI22M1P U201 ( .A(\Queue[1][10] ), .B(n92), .C(n5), .D(Packet_Out[10]), .Z(
        n70) );
  OAI21M1P U202 ( .A(n161), .B(n94), .C(n70), .Z(n452) );
  AOI22M1P U203 ( .A(\Queue[1][11] ), .B(n92), .C(n91), .D(Packet_Out[11]), 
        .Z(n71) );
  OAI21M1P U204 ( .A(n163), .B(n94), .C(n71), .Z(n453) );
  AOI22M1P U205 ( .A(\Queue[1][12] ), .B(n92), .C(n91), .D(Packet_Out[12]), 
        .Z(n72) );
  OAI21M1P U206 ( .A(n165), .B(n94), .C(n72), .Z(n454) );
  AOI22M1P U207 ( .A(\Queue[1][13] ), .B(n92), .C(n91), .D(Packet_Out[13]), 
        .Z(n73) );
  OAI21M1P U208 ( .A(n167), .B(n94), .C(n73), .Z(n455) );
  AOI22M1P U209 ( .A(\Queue[1][14] ), .B(n92), .C(n91), .D(Packet_Out[14]), 
        .Z(n74) );
  OAI21M1P U210 ( .A(n169), .B(n94), .C(n74), .Z(n456) );
  AOI22M1P U211 ( .A(\Queue[1][15] ), .B(n92), .C(n91), .D(Packet_Out[15]), 
        .Z(n75) );
  OAI21M1P U212 ( .A(n171), .B(n94), .C(n75), .Z(n457) );
  AOI22M1P U213 ( .A(\Queue[1][16] ), .B(n92), .C(n91), .D(Packet_Out[16]), 
        .Z(n76) );
  OAI21M1P U214 ( .A(n173), .B(n94), .C(n76), .Z(n458) );
  AOI22M1P U215 ( .A(\Queue[1][17] ), .B(n92), .C(n91), .D(Packet_Out[17]), 
        .Z(n77) );
  OAI21M1P U216 ( .A(n175), .B(n94), .C(n77), .Z(n459) );
  AOI22M1P U217 ( .A(\Queue[1][18] ), .B(n92), .C(n91), .D(Packet_Out[18]), 
        .Z(n78) );
  OAI21M1P U218 ( .A(n177), .B(n94), .C(n78), .Z(n460) );
  AOI22M1P U219 ( .A(\Queue[1][19] ), .B(n92), .C(n91), .D(Packet_Out[19]), 
        .Z(n79) );
  OAI21M1P U220 ( .A(n179), .B(n94), .C(n79), .Z(n461) );
  AOI22M1P U221 ( .A(\Queue[1][20] ), .B(n92), .C(n5), .D(Packet_Out[20]), .Z(
        n80) );
  OAI21M1P U222 ( .A(n181), .B(n94), .C(n80), .Z(n462) );
  AOI22M1P U223 ( .A(\Queue[1][21] ), .B(n92), .C(n5), .D(Packet_Out[21]), .Z(
        n81) );
  OAI21M1P U224 ( .A(n183), .B(n94), .C(n81), .Z(n463) );
  AOI22M1P U225 ( .A(\Queue[1][22] ), .B(n92), .C(n5), .D(Packet_Out[22]), .Z(
        n82) );
  OAI21M1P U226 ( .A(n185), .B(n94), .C(n82), .Z(n464) );
  AOI22M1P U227 ( .A(\Queue[1][23] ), .B(n92), .C(n5), .D(Packet_Out[23]), .Z(
        n83) );
  OAI21M1P U228 ( .A(n187), .B(n94), .C(n83), .Z(n465) );
  AOI22M1P U229 ( .A(\Queue[1][24] ), .B(n92), .C(n5), .D(Packet_Out[24]), .Z(
        n84) );
  OAI21M1P U230 ( .A(n189), .B(n94), .C(n84), .Z(n466) );
  AOI22M1P U231 ( .A(\Queue[1][25] ), .B(n92), .C(n5), .D(Packet_Out[25]), .Z(
        n85) );
  OAI21M1P U232 ( .A(n191), .B(n94), .C(n85), .Z(n467) );
  AOI22M1P U233 ( .A(\Queue[1][26] ), .B(n92), .C(n5), .D(Packet_Out[26]), .Z(
        n86) );
  OAI21M1P U234 ( .A(n193), .B(n94), .C(n86), .Z(n468) );
  AOI22M1P U235 ( .A(\Queue[1][27] ), .B(n92), .C(n5), .D(Packet_Out[27]), .Z(
        n87) );
  OAI21M1P U236 ( .A(n195), .B(n94), .C(n87), .Z(n469) );
  AOI22M1P U237 ( .A(\Queue[1][28] ), .B(n92), .C(n5), .D(Packet_Out[28]), .Z(
        n88) );
  OAI21M1P U238 ( .A(n197), .B(n94), .C(n88), .Z(n470) );
  AOI22M1P U239 ( .A(\Queue[1][29] ), .B(n92), .C(n5), .D(Packet_Out[29]), .Z(
        n89) );
  OAI21M1P U240 ( .A(n199), .B(n94), .C(n89), .Z(n471) );
  AOI22M1P U241 ( .A(\Queue[1][30] ), .B(n92), .C(n91), .D(Packet_Out[30]), 
        .Z(n90) );
  OAI21M1P U242 ( .A(n201), .B(n94), .C(n90), .Z(n472) );
  AOI22M1P U243 ( .A(\Queue[1][31] ), .B(n92), .C(n5), .D(Packet_Out[31]), .Z(
        n93) );
  OAI21M1P U244 ( .A(n206), .B(n94), .C(n93), .Z(n473) );
  OA21M1P U245 ( .A(n136), .B(n97), .C(Rst_n), .Z(n95) );
  ND2M1P U246 ( .A(n96), .B(n134), .Z(n135) );
  AOI22M1P U247 ( .A(\Queue[2][0] ), .B(n6), .C(\Queue[3][0] ), .D(n129), .Z(
        n98) );
  OAI21M1P U248 ( .A(n141), .B(n132), .C(n98), .Z(n474) );
  OAI21M1P U249 ( .A(n143), .B(n132), .C(n99), .Z(n475) );
  AOI22M1P U250 ( .A(\Queue[2][2] ), .B(n6), .C(n129), .D(\Queue[3][2] ), .Z(
        n100) );
  OAI21M1P U251 ( .A(n145), .B(n132), .C(n100), .Z(n476) );
  AOI22M1P U252 ( .A(\Queue[2][3] ), .B(n6), .C(n129), .D(\Queue[3][3] ), .Z(
        n101) );
  OAI21M1P U253 ( .A(n147), .B(n132), .C(n101), .Z(n477) );
  AOI22M1P U254 ( .A(\Queue[2][4] ), .B(n6), .C(n129), .D(\Queue[3][4] ), .Z(
        n102) );
  OAI21M1P U255 ( .A(n149), .B(n132), .C(n102), .Z(n478) );
  AOI22M1P U256 ( .A(\Queue[2][5] ), .B(n6), .C(n129), .D(\Queue[3][5] ), .Z(
        n103) );
  OAI21M1P U257 ( .A(n151), .B(n132), .C(n103), .Z(n479) );
  AOI22M1P U258 ( .A(\Queue[2][6] ), .B(n6), .C(n129), .D(\Queue[3][6] ), .Z(
        n104) );
  OAI21M1P U259 ( .A(n153), .B(n132), .C(n104), .Z(n480) );
  AOI22M1P U260 ( .A(\Queue[2][7] ), .B(n6), .C(n129), .D(\Queue[3][7] ), .Z(
        n105) );
  OAI21M1P U261 ( .A(n155), .B(n132), .C(n105), .Z(n481) );
  AOI22M1P U262 ( .A(\Queue[2][8] ), .B(n6), .C(n129), .D(\Queue[3][8] ), .Z(
        n106) );
  OAI21M1P U263 ( .A(n157), .B(n132), .C(n106), .Z(n482) );
  AOI22M1P U264 ( .A(\Queue[2][9] ), .B(n6), .C(n129), .D(\Queue[3][9] ), .Z(
        n107) );
  OAI21M1P U265 ( .A(n159), .B(n132), .C(n107), .Z(n483) );
  AOI22M1P U266 ( .A(\Queue[2][10] ), .B(n6), .C(n129), .D(\Queue[3][10] ), 
        .Z(n108) );
  OAI21M1P U267 ( .A(n161), .B(n132), .C(n108), .Z(n484) );
  AOI22M1P U268 ( .A(\Queue[2][11] ), .B(n6), .C(n129), .D(\Queue[3][11] ), 
        .Z(n109) );
  OAI21M1P U269 ( .A(n163), .B(n132), .C(n109), .Z(n485) );
  AOI22M1P U270 ( .A(\Queue[2][12] ), .B(n6), .C(n129), .D(\Queue[3][12] ), 
        .Z(n110) );
  OAI21M1P U271 ( .A(n165), .B(n132), .C(n110), .Z(n486) );
  AOI22M1P U272 ( .A(\Queue[2][13] ), .B(n6), .C(n129), .D(\Queue[3][13] ), 
        .Z(n111) );
  OAI21M1P U273 ( .A(n167), .B(n132), .C(n111), .Z(n487) );
  AOI22M1P U274 ( .A(\Queue[2][14] ), .B(n6), .C(n129), .D(\Queue[3][14] ), 
        .Z(n112) );
  OAI21M1P U275 ( .A(n169), .B(n132), .C(n112), .Z(n488) );
  AOI22M1P U276 ( .A(\Queue[2][15] ), .B(n6), .C(n129), .D(\Queue[3][15] ), 
        .Z(n113) );
  OAI21M1P U277 ( .A(n171), .B(n132), .C(n113), .Z(n489) );
  AOI22M1P U278 ( .A(\Queue[2][16] ), .B(n6), .C(n129), .D(\Queue[3][16] ), 
        .Z(n114) );
  OAI21M1P U279 ( .A(n173), .B(n132), .C(n114), .Z(n490) );
  AOI22M1P U280 ( .A(\Queue[2][17] ), .B(n6), .C(n129), .D(\Queue[3][17] ), 
        .Z(n115) );
  OAI21M1P U281 ( .A(n175), .B(n132), .C(n115), .Z(n491) );
  AOI22M1P U282 ( .A(\Queue[2][18] ), .B(n6), .C(n129), .D(\Queue[3][18] ), 
        .Z(n116) );
  OAI21M1P U283 ( .A(n177), .B(n132), .C(n116), .Z(n492) );
  AOI22M1P U284 ( .A(\Queue[2][19] ), .B(n6), .C(n129), .D(\Queue[3][19] ), 
        .Z(n117) );
  OAI21M1P U285 ( .A(n179), .B(n132), .C(n117), .Z(n493) );
  AOI22M1P U286 ( .A(\Queue[2][20] ), .B(n7), .C(n129), .D(\Queue[3][20] ), 
        .Z(n118) );
  OAI21M1P U287 ( .A(n181), .B(n132), .C(n118), .Z(n494) );
  AOI22M1P U288 ( .A(\Queue[2][21] ), .B(n7), .C(n129), .D(\Queue[3][21] ), 
        .Z(n119) );
  OAI21M1P U289 ( .A(n183), .B(n132), .C(n119), .Z(n495) );
  AOI22M1P U290 ( .A(\Queue[2][22] ), .B(n7), .C(n129), .D(\Queue[3][22] ), 
        .Z(n120) );
  OAI21M1P U291 ( .A(n185), .B(n132), .C(n120), .Z(n496) );
  AOI22M1P U292 ( .A(\Queue[2][23] ), .B(n7), .C(n129), .D(\Queue[3][23] ), 
        .Z(n121) );
  OAI21M1P U293 ( .A(n187), .B(n132), .C(n121), .Z(n497) );
  AOI22M1P U294 ( .A(\Queue[2][24] ), .B(n7), .C(n129), .D(\Queue[3][24] ), 
        .Z(n122) );
  OAI21M1P U295 ( .A(n189), .B(n132), .C(n122), .Z(n498) );
  AOI22M1P U296 ( .A(\Queue[2][25] ), .B(n7), .C(n129), .D(\Queue[3][25] ), 
        .Z(n123) );
  OAI21M1P U297 ( .A(n191), .B(n132), .C(n123), .Z(n499) );
  AOI22M1P U298 ( .A(\Queue[2][26] ), .B(n7), .C(n129), .D(\Queue[3][26] ), 
        .Z(n124) );
  OAI21M1P U299 ( .A(n193), .B(n132), .C(n124), .Z(n500) );
  AOI22M1P U300 ( .A(\Queue[2][27] ), .B(n7), .C(n129), .D(\Queue[3][27] ), 
        .Z(n125) );
  OAI21M1P U301 ( .A(n195), .B(n132), .C(n125), .Z(n501) );
  AOI22M1P U302 ( .A(\Queue[2][28] ), .B(n7), .C(n129), .D(\Queue[3][28] ), 
        .Z(n126) );
  OAI21M1P U303 ( .A(n197), .B(n132), .C(n126), .Z(n502) );
  AOI22M1P U304 ( .A(\Queue[2][29] ), .B(n7), .C(n129), .D(\Queue[3][29] ), 
        .Z(n127) );
  OAI21M1P U305 ( .A(n199), .B(n132), .C(n127), .Z(n503) );
  AOI22M1P U306 ( .A(\Queue[2][30] ), .B(n6), .C(n129), .D(\Queue[3][30] ), 
        .Z(n128) );
  OAI21M1P U307 ( .A(n201), .B(n132), .C(n128), .Z(n504) );
  AOI22M1P U308 ( .A(\Queue[2][31] ), .B(n7), .C(n129), .D(\Queue[3][31] ), 
        .Z(n131) );
  OAI21M1P U309 ( .A(n206), .B(n132), .C(n131), .Z(n505) );
  OA21M1P U310 ( .A(n136), .B(n137), .C(Rst_n), .Z(n133) );
  AOI22M1P U311 ( .A(\Queue[3][0] ), .B(n8), .C(n202), .D(\Queue[4][0] ), .Z(
        n140) );
  OAI21M1P U312 ( .A(n141), .B(n205), .C(n140), .Z(n506) );
  AOI22M1P U313 ( .A(\Queue[3][1] ), .B(n8), .C(n202), .D(\Queue[4][1] ), .Z(
        n142) );
  OAI21M1P U314 ( .A(n143), .B(n205), .C(n142), .Z(n507) );
  AOI22M1P U315 ( .A(\Queue[3][2] ), .B(n8), .C(n202), .D(\Queue[4][2] ), .Z(
        n144) );
  OAI21M1P U316 ( .A(n145), .B(n205), .C(n144), .Z(n508) );
  AOI22M1P U317 ( .A(\Queue[3][3] ), .B(n8), .C(n202), .D(\Queue[4][3] ), .Z(
        n146) );
  OAI21M1P U318 ( .A(n147), .B(n205), .C(n146), .Z(n509) );
  AOI22M1P U319 ( .A(\Queue[3][4] ), .B(n8), .C(n202), .D(\Queue[4][4] ), .Z(
        n148) );
  OAI21M1P U320 ( .A(n149), .B(n205), .C(n148), .Z(n510) );
  AOI22M1P U321 ( .A(\Queue[3][5] ), .B(n8), .C(n202), .D(\Queue[4][5] ), .Z(
        n150) );
  OAI21M1P U322 ( .A(n151), .B(n205), .C(n150), .Z(n511) );
  AOI22M1P U323 ( .A(\Queue[3][6] ), .B(n8), .C(n202), .D(\Queue[4][6] ), .Z(
        n152) );
  OAI21M1P U324 ( .A(n153), .B(n205), .C(n152), .Z(n512) );
  AOI22M1P U325 ( .A(\Queue[3][7] ), .B(n8), .C(n202), .D(\Queue[4][7] ), .Z(
        n154) );
  OAI21M1P U326 ( .A(n155), .B(n205), .C(n154), .Z(n513) );
  AOI22M1P U327 ( .A(\Queue[3][8] ), .B(n8), .C(n202), .D(\Queue[4][8] ), .Z(
        n156) );
  OAI21M1P U328 ( .A(n157), .B(n205), .C(n156), .Z(n514) );
  AOI22M1P U329 ( .A(\Queue[3][9] ), .B(n8), .C(n202), .D(\Queue[4][9] ), .Z(
        n158) );
  OAI21M1P U330 ( .A(n159), .B(n205), .C(n158), .Z(n515) );
  AOI22M1P U331 ( .A(\Queue[3][10] ), .B(n8), .C(n202), .D(\Queue[4][10] ), 
        .Z(n160) );
  OAI21M1P U332 ( .A(n161), .B(n205), .C(n160), .Z(n516) );
  AOI22M1P U333 ( .A(\Queue[3][11] ), .B(n8), .C(n202), .D(\Queue[4][11] ), 
        .Z(n162) );
  OAI21M1P U334 ( .A(n163), .B(n205), .C(n162), .Z(n517) );
  AOI22M1P U335 ( .A(\Queue[3][12] ), .B(n8), .C(n202), .D(\Queue[4][12] ), 
        .Z(n164) );
  OAI21M1P U336 ( .A(n165), .B(n205), .C(n164), .Z(n518) );
  AOI22M1P U337 ( .A(\Queue[3][13] ), .B(n8), .C(n202), .D(\Queue[4][13] ), 
        .Z(n166) );
  OAI21M1P U338 ( .A(n167), .B(n205), .C(n166), .Z(n519) );
  AOI22M1P U339 ( .A(\Queue[3][14] ), .B(n8), .C(n202), .D(\Queue[4][14] ), 
        .Z(n168) );
  OAI21M1P U340 ( .A(n169), .B(n205), .C(n168), .Z(n520) );
  AOI22M1P U341 ( .A(\Queue[3][15] ), .B(n8), .C(n202), .D(\Queue[4][15] ), 
        .Z(n170) );
  OAI21M1P U342 ( .A(n171), .B(n205), .C(n170), .Z(n521) );
  AOI22M1P U343 ( .A(\Queue[3][16] ), .B(n8), .C(n202), .D(\Queue[4][16] ), 
        .Z(n172) );
  OAI21M1P U344 ( .A(n173), .B(n205), .C(n172), .Z(n522) );
  AOI22M1P U345 ( .A(\Queue[3][17] ), .B(n8), .C(n202), .D(\Queue[4][17] ), 
        .Z(n174) );
  OAI21M1P U346 ( .A(n175), .B(n205), .C(n174), .Z(n523) );
  AOI22M1P U347 ( .A(\Queue[3][18] ), .B(n8), .C(n202), .D(\Queue[4][18] ), 
        .Z(n176) );
  OAI21M1P U348 ( .A(n177), .B(n205), .C(n176), .Z(n524) );
  AOI22M1P U349 ( .A(\Queue[3][19] ), .B(n8), .C(n202), .D(\Queue[4][19] ), 
        .Z(n178) );
  OAI21M1P U350 ( .A(n179), .B(n205), .C(n178), .Z(n525) );
  AOI22M1P U351 ( .A(\Queue[3][20] ), .B(n9), .C(n202), .D(\Queue[4][20] ), 
        .Z(n180) );
  OAI21M1P U352 ( .A(n181), .B(n205), .C(n180), .Z(n526) );
  AOI22M1P U353 ( .A(\Queue[3][21] ), .B(n9), .C(n202), .D(\Queue[4][21] ), 
        .Z(n182) );
  OAI21M1P U354 ( .A(n183), .B(n205), .C(n182), .Z(n527) );
  AOI22M1P U355 ( .A(\Queue[3][22] ), .B(n9), .C(n202), .D(\Queue[4][22] ), 
        .Z(n184) );
  OAI21M1P U356 ( .A(n185), .B(n205), .C(n184), .Z(n528) );
  AOI22M1P U357 ( .A(\Queue[3][23] ), .B(n9), .C(n202), .D(\Queue[4][23] ), 
        .Z(n186) );
  OAI21M1P U358 ( .A(n187), .B(n205), .C(n186), .Z(n529) );
  AOI22M1P U359 ( .A(\Queue[3][24] ), .B(n9), .C(n202), .D(\Queue[4][24] ), 
        .Z(n188) );
  OAI21M1P U360 ( .A(n189), .B(n205), .C(n188), .Z(n530) );
  AOI22M1P U361 ( .A(\Queue[3][25] ), .B(n9), .C(n202), .D(\Queue[4][25] ), 
        .Z(n190) );
  OAI21M1P U362 ( .A(n191), .B(n205), .C(n190), .Z(n531) );
  AOI22M1P U363 ( .A(\Queue[3][26] ), .B(n9), .C(n202), .D(\Queue[4][26] ), 
        .Z(n192) );
  OAI21M1P U364 ( .A(n193), .B(n205), .C(n192), .Z(n532) );
  AOI22M1P U365 ( .A(\Queue[3][27] ), .B(n9), .C(n202), .D(\Queue[4][27] ), 
        .Z(n194) );
  OAI21M1P U366 ( .A(n195), .B(n205), .C(n194), .Z(n533) );
  AOI22M1P U367 ( .A(\Queue[3][28] ), .B(n9), .C(n202), .D(\Queue[4][28] ), 
        .Z(n196) );
  OAI21M1P U368 ( .A(n197), .B(n205), .C(n196), .Z(n534) );
  AOI22M1P U369 ( .A(\Queue[3][29] ), .B(n9), .C(n202), .D(\Queue[4][29] ), 
        .Z(n198) );
  OAI21M1P U370 ( .A(n199), .B(n205), .C(n198), .Z(n535) );
  AOI22M1P U371 ( .A(\Queue[3][30] ), .B(n8), .C(n202), .D(\Queue[4][30] ), 
        .Z(n200) );
  OAI21M1P U372 ( .A(n201), .B(n205), .C(n200), .Z(n536) );
  AOI22M1P U373 ( .A(\Queue[3][31] ), .B(n9), .C(n202), .D(\Queue[4][31] ), 
        .Z(n204) );
  OAI21M1P U374 ( .A(n206), .B(n205), .C(n204), .Z(n537) );
  AOI22M1P U375 ( .A(n373), .B(n208), .C(n207), .D(Empty), .Z(n539) );
endmodule


module Link_Control_0 ( Clk_r, Rst_n, Tx_Ready, Tx_Error, RxData_Valid, RxData, 
        Packet_From_Core, TxQueue_Write, RxQueue_Read, TxData_Valid, TxData, 
        Error_Ack, Core_Rcv_Ready, Packet_To_Core, RxQueue_Empty, TxQueue_Full
 );
  input [31:0] RxData;
  input [31:0] Packet_From_Core;
  output [31:0] TxData;
  output [31:0] Packet_To_Core;
  input Clk_r, Rst_n, Tx_Ready, Tx_Error, RxData_Valid, TxQueue_Write,
         RxQueue_Read;
  output TxData_Valid, Error_Ack, Core_Rcv_Ready, RxQueue_Empty, TxQueue_Full;
  wire   TxQueue_Read, TxQueue_Empty, RxQueue_Write, RxQueue_Full, N9, N16, n1,
         n2, n3, n4, n5;

  Packet_Queue_0 TxQueue ( .Clk_r(Clk_r), .Rst_n(Rst_n), .Packet_In(
        Packet_From_Core), .Read_Ack(TxQueue_Read), .Write_Ack(TxQueue_Write), 
        .Packet_Out(TxData), .Empty(TxQueue_Empty), .Full(TxQueue_Full) );
  Packet_Queue_9 RxQueue ( .Clk_r(Clk_r), .Rst_n(Rst_n), .Packet_In(RxData), 
        .Read_Ack(RxQueue_Read), .Write_Ack(RxQueue_Write), .Packet_Out(
        Packet_To_Core), .Empty(RxQueue_Empty), .Full(RxQueue_Full) );
  FD4QM1P TxData_Valid_reg ( .D(n1), .CP(Clk_r), .SD(Rst_n), .Q(n2) );
  FD4QM1P RxQueue_Write_reg ( .D(n3), .CP(Clk_r), .SD(Rst_n), .Q(n4) );
  FD2QM1P TxQueue_Read_reg ( .D(N16), .CP(Clk_r), .CD(Rst_n), .Q(TxQueue_Read)
         );
  FD2QM1P Core_Rcv_Ready_reg ( .D(N9), .CP(Clk_r), .CD(Rst_n), .Q(
        Core_Rcv_Ready) );
  N1M4P U3 ( .A(n4), .Z(RxQueue_Write) );
  NR2M1P U4 ( .A(n2), .B(Tx_Ready), .Z(N16) );
  NR2M1P U5 ( .A(RxData_Valid), .B(RxQueue_Full), .Z(n5) );
  OA21M1P U6 ( .A(Core_Rcv_Ready), .B(n5), .C(n4), .Z(N9) );
  N1M1P U7 ( .A(n2), .Z(TxData_Valid) );
  ND3M1P U8 ( .A(n4), .B(Core_Rcv_Ready), .C(RxData_Valid), .Z(n3) );
  AO21CNM1P U9 ( .A(n2), .B(TxQueue_Empty), .C(Tx_Ready), .Z(n1) );
endmodule


module Routing_State_Machine ( Clk_r, Rst_n, Router_Address, Link_Config, 
        Packet_From_Link_N, Packet_From_Link_S, Packet_From_Link_W, 
        Packet_From_Link_E, Packet_From_Node, RxQueue_Empty_N, RxQueue_Empty_S, 
        RxQueue_Empty_W, RxQueue_Empty_E, TxQueue_Full_N, TxQueue_Full_S, 
        TxQueue_Full_W, TxQueue_Full_E, To_Node_Full, Node_Queue_Empty, 
        Packet_To_Link_N, Packet_To_Link_S, Packet_To_Link_W, Packet_To_Link_E, 
        Packet_To_Node, TxQueue_Write_N, TxQueue_Write_S, TxQueue_Write_W, 
        TxQueue_Write_E, To_Node_Write, RxQueue_Read_N, RxQueue_Read_S, 
        RxQueue_Read_W, RxQueue_Read_E, Node_Read );
  input [7:0] Router_Address;
  input [3:0] Link_Config;
  input [31:0] Packet_From_Link_N;
  input [31:0] Packet_From_Link_S;
  input [31:0] Packet_From_Link_W;
  input [31:0] Packet_From_Link_E;
  input [31:0] Packet_From_Node;
  output [31:0] Packet_To_Link_N;
  output [31:0] Packet_To_Link_S;
  output [31:0] Packet_To_Link_W;
  output [31:0] Packet_To_Link_E;
  output [31:0] Packet_To_Node;
  input Clk_r, Rst_n, RxQueue_Empty_N, RxQueue_Empty_S, RxQueue_Empty_W,
         RxQueue_Empty_E, TxQueue_Full_N, TxQueue_Full_S, TxQueue_Full_W,
         TxQueue_Full_E, To_Node_Full, Node_Queue_Empty;
  output TxQueue_Write_N, TxQueue_Write_S, TxQueue_Write_W, TxQueue_Write_E,
         To_Node_Write, RxQueue_Read_N, RxQueue_Read_S, RxQueue_Read_W,
         RxQueue_Read_E, Node_Read;
  wire   Packet_From_Node_31, Packet_From_Node_30, Packet_From_Node_29,
         Packet_From_Node_28, Packet_From_Node_27, Packet_From_Node_26,
         Packet_From_Node_25, Packet_From_Node_24, N43, N44, N48, N108, N109,
         N110, N111, N112, N113, N114, N115, n1, n2, n3, n4, n5, n6, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n32, n33, n34, n35, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n57, n107, n245, n246, n247, n249,
         n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
         n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n31, n36, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n248, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307;
  wire   [31:0] chosenPacket;
  wire   [2:0] dataLocation;
  assign Packet_From_Node_31 = Packet_From_Node[31];
  assign Packet_From_Node_30 = Packet_From_Node[30];
  assign Packet_From_Node_29 = Packet_From_Node[29];
  assign Packet_From_Node_28 = Packet_From_Node[28];
  assign Packet_From_Node_27 = Packet_From_Node[27];
  assign Packet_From_Node_26 = Packet_From_Node[26];
  assign Packet_From_Node_25 = Packet_From_Node[25];
  assign Packet_From_Node_24 = Packet_From_Node[24];

  FD2LQM1P \dataLocation_reg[0]  ( .D(N43), .LD(n8), .CP(Clk_r), .CD(Rst_n), 
        .Q(dataLocation[0]) );
  FD4QM1P \Packet_To_Node_reg[16]  ( .D(n25), .CP(Clk_r), .SD(Rst_n), .Q(
        Packet_To_Node[16]) );
  FD4QM1P \Packet_To_Node_reg[17]  ( .D(n26), .CP(Clk_r), .SD(Rst_n), .Q(
        Packet_To_Node[17]) );
  FD4QM1P \Packet_To_Node_reg[18]  ( .D(n27), .CP(Clk_r), .SD(Rst_n), .Q(
        Packet_To_Node[18]) );
  FD4QM1P \Packet_To_Node_reg[19]  ( .D(n28), .CP(Clk_r), .SD(Rst_n), .Q(
        Packet_To_Node[19]) );
  FD4QM1P \Packet_To_Node_reg[20]  ( .D(n29), .CP(Clk_r), .SD(Rst_n), .Q(
        Packet_To_Node[20]) );
  FD4QM1P \Packet_To_Node_reg[21]  ( .D(n30), .CP(Clk_r), .SD(Rst_n), .Q(
        Packet_To_Node[21]) );
  FD4QM1P \Packet_To_Node_reg[23]  ( .D(n32), .CP(Clk_r), .SD(Rst_n), .Q(
        Packet_To_Node[23]) );
  FD2LQM1P \dataLocation_reg[1]  ( .D(N44), .LD(n8), .CP(Clk_r), .CD(Rst_n), 
        .Q(dataLocation[1]) );
  FD2LQM1P \dataLocation_reg[2]  ( .D(n57), .LD(n8), .CP(Clk_r), .CD(Rst_n), 
        .Q(n6) );
  FD1QM1P \chosenPacket_reg[31]  ( .D(n263), .CP(Clk_r), .Q(chosenPacket[31])
         );
  FD2LQM1P \Packet_To_Node_reg[31]  ( .D(n41), .LD(n65), .CP(Clk_r), .CD(Rst_n), .Q(n5) );
  FD1QM1P \chosenPacket_reg[30]  ( .D(n264), .CP(Clk_r), .Q(chosenPacket[30])
         );
  FD2LQM1P \Packet_To_Node_reg[30]  ( .D(n42), .LD(n65), .CP(Clk_r), .CD(Rst_n), .Q(n4) );
  FD1QM1P \chosenPacket_reg[29]  ( .D(n265), .CP(Clk_r), .Q(chosenPacket[29])
         );
  FD2LQM1P \Packet_To_Node_reg[29]  ( .D(n43), .LD(n65), .CP(Clk_r), .CD(Rst_n), .Q(n3) );
  FD1QM1P \chosenPacket_reg[28]  ( .D(n266), .CP(Clk_r), .Q(chosenPacket[28])
         );
  FD4QM1P \Packet_To_Node_reg[28]  ( .D(n35), .CP(Clk_r), .SD(Rst_n), .Q(
        Packet_To_Node[28]) );
  FD1QM1P \chosenPacket_reg[27]  ( .D(n267), .CP(Clk_r), .Q(chosenPacket[27])
         );
  FD2LQM1P \Packet_To_Node_reg[27]  ( .D(n44), .LD(n65), .CP(Clk_r), .CD(Rst_n), .Q(n2) );
  FD1QM1P \chosenPacket_reg[26]  ( .D(n268), .CP(Clk_r), .Q(chosenPacket[26])
         );
  FD4QM1P \Packet_To_Node_reg[26]  ( .D(n34), .CP(Clk_r), .SD(Rst_n), .Q(
        Packet_To_Node[26]) );
  FD1QM1P \chosenPacket_reg[25]  ( .D(n269), .CP(Clk_r), .Q(chosenPacket[25])
         );
  FD2LQM1P \Packet_To_Node_reg[25]  ( .D(n45), .LD(n65), .CP(Clk_r), .CD(Rst_n), .Q(n1) );
  FD1QM1P \chosenPacket_reg[24]  ( .D(n270), .CP(Clk_r), .Q(chosenPacket[24])
         );
  FD1LQM1P \Packet_To_Link_N_reg[31]  ( .D(chosenPacket[31]), .LD(n39), .CP(
        Clk_r), .Q(Packet_To_Link_N[31]) );
  FD1LQM1P \Packet_To_Link_N_reg[30]  ( .D(chosenPacket[30]), .LD(n39), .CP(
        Clk_r), .Q(Packet_To_Link_N[30]) );
  FD1LQM1P \Packet_To_Link_N_reg[29]  ( .D(chosenPacket[29]), .LD(n39), .CP(
        Clk_r), .Q(Packet_To_Link_N[29]) );
  FD1LQM1P \Packet_To_Link_N_reg[27]  ( .D(chosenPacket[27]), .LD(n39), .CP(
        Clk_r), .Q(Packet_To_Link_N[27]) );
  FD1LQM1P \Packet_To_Link_N_reg[25]  ( .D(chosenPacket[25]), .LD(n39), .CP(
        Clk_r), .Q(Packet_To_Link_N[25]) );
  FD1LQM1P \Packet_To_Link_N_reg[16]  ( .D(N108), .LD(n39), .CP(Clk_r), .Q(
        Packet_To_Link_N[16]) );
  FD1LQM1P \Packet_To_Link_N_reg[17]  ( .D(N109), .LD(n39), .CP(Clk_r), .Q(
        Packet_To_Link_N[17]) );
  FD1LQM1P \Packet_To_Link_N_reg[18]  ( .D(N110), .LD(n39), .CP(Clk_r), .Q(
        Packet_To_Link_N[18]) );
  FD1LQM1P \Packet_To_Link_N_reg[19]  ( .D(N111), .LD(n39), .CP(Clk_r), .Q(
        Packet_To_Link_N[19]) );
  FD1LQM1P \Packet_To_Link_N_reg[20]  ( .D(N112), .LD(n39), .CP(Clk_r), .Q(
        Packet_To_Link_N[20]) );
  FD1LQM1P \Packet_To_Link_N_reg[21]  ( .D(N113), .LD(n39), .CP(Clk_r), .Q(
        Packet_To_Link_N[21]) );
  FD1LQM1P \Packet_To_Link_N_reg[22]  ( .D(N114), .LD(n39), .CP(Clk_r), .Q(
        Packet_To_Link_N[22]) );
  FD1LQM1P \Packet_To_Link_N_reg[23]  ( .D(N115), .LD(n39), .CP(Clk_r), .Q(
        Packet_To_Link_N[23]) );
  FD1LQM1P \Packet_To_Link_N_reg[26]  ( .D(chosenPacket[26]), .LD(n39), .CP(
        Clk_r), .Q(Packet_To_Link_N[26]) );
  FD1LQM1P \Packet_To_Link_N_reg[28]  ( .D(chosenPacket[28]), .LD(n39), .CP(
        Clk_r), .Q(Packet_To_Link_N[28]) );
  FD1LQM1P \Packet_To_Link_S_reg[31]  ( .D(chosenPacket[31]), .LD(n40), .CP(
        Clk_r), .Q(Packet_To_Link_S[31]) );
  FD1LQM1P \Packet_To_Link_S_reg[30]  ( .D(chosenPacket[30]), .LD(n40), .CP(
        Clk_r), .Q(Packet_To_Link_S[30]) );
  FD1LQM1P \Packet_To_Link_S_reg[29]  ( .D(chosenPacket[29]), .LD(n40), .CP(
        Clk_r), .Q(Packet_To_Link_S[29]) );
  FD1LQM1P \Packet_To_Link_S_reg[27]  ( .D(chosenPacket[27]), .LD(n40), .CP(
        Clk_r), .Q(Packet_To_Link_S[27]) );
  FD1LQM1P \Packet_To_Link_S_reg[25]  ( .D(chosenPacket[25]), .LD(n40), .CP(
        Clk_r), .Q(Packet_To_Link_S[25]) );
  FD1LQM1P \Packet_To_Link_S_reg[16]  ( .D(N108), .LD(n40), .CP(Clk_r), .Q(
        Packet_To_Link_S[16]) );
  FD1LQM1P \Packet_To_Link_S_reg[17]  ( .D(N109), .LD(n40), .CP(Clk_r), .Q(
        Packet_To_Link_S[17]) );
  FD1LQM1P \Packet_To_Link_S_reg[18]  ( .D(N110), .LD(n40), .CP(Clk_r), .Q(
        Packet_To_Link_S[18]) );
  FD1LQM1P \Packet_To_Link_S_reg[19]  ( .D(N111), .LD(n40), .CP(Clk_r), .Q(
        Packet_To_Link_S[19]) );
  FD1LQM1P \Packet_To_Link_S_reg[20]  ( .D(N112), .LD(n40), .CP(Clk_r), .Q(
        Packet_To_Link_S[20]) );
  FD1LQM1P \Packet_To_Link_S_reg[21]  ( .D(N113), .LD(n40), .CP(Clk_r), .Q(
        Packet_To_Link_S[21]) );
  FD1LQM1P \Packet_To_Link_S_reg[22]  ( .D(N114), .LD(n40), .CP(Clk_r), .Q(
        Packet_To_Link_S[22]) );
  FD1LQM1P \Packet_To_Link_S_reg[23]  ( .D(N115), .LD(n40), .CP(Clk_r), .Q(
        Packet_To_Link_S[23]) );
  FD1LQM1P \Packet_To_Link_S_reg[26]  ( .D(chosenPacket[26]), .LD(n40), .CP(
        Clk_r), .Q(Packet_To_Link_S[26]) );
  FD1LQM1P \Packet_To_Link_S_reg[28]  ( .D(chosenPacket[28]), .LD(n40), .CP(
        Clk_r), .Q(Packet_To_Link_S[28]) );
  FD1LQM1P \Packet_To_Link_W_reg[31]  ( .D(chosenPacket[31]), .LD(n68), .CP(
        Clk_r), .Q(Packet_To_Link_W[31]) );
  FD1LQM1P \Packet_To_Link_W_reg[30]  ( .D(chosenPacket[30]), .LD(n67), .CP(
        Clk_r), .Q(Packet_To_Link_W[30]) );
  FD1LQM1P \Packet_To_Link_W_reg[29]  ( .D(chosenPacket[29]), .LD(n68), .CP(
        Clk_r), .Q(Packet_To_Link_W[29]) );
  FD1LQM1P \Packet_To_Link_W_reg[27]  ( .D(chosenPacket[27]), .LD(n67), .CP(
        Clk_r), .Q(Packet_To_Link_W[27]) );
  FD1LQM1P \Packet_To_Link_W_reg[25]  ( .D(chosenPacket[25]), .LD(n68), .CP(
        Clk_r), .Q(Packet_To_Link_W[25]) );
  FD1LQM1P \Packet_To_Link_W_reg[16]  ( .D(N108), .LD(n67), .CP(Clk_r), .Q(
        Packet_To_Link_W[16]) );
  FD1LQM1P \Packet_To_Link_W_reg[17]  ( .D(N109), .LD(n68), .CP(Clk_r), .Q(
        Packet_To_Link_W[17]) );
  FD1LQM1P \Packet_To_Link_W_reg[18]  ( .D(N110), .LD(n67), .CP(Clk_r), .Q(
        Packet_To_Link_W[18]) );
  FD1LQM1P \Packet_To_Link_W_reg[19]  ( .D(N111), .LD(n68), .CP(Clk_r), .Q(
        Packet_To_Link_W[19]) );
  FD1LQM1P \Packet_To_Link_W_reg[20]  ( .D(N112), .LD(n67), .CP(Clk_r), .Q(
        Packet_To_Link_W[20]) );
  FD1LQM1P \Packet_To_Link_W_reg[21]  ( .D(N113), .LD(n68), .CP(Clk_r), .Q(
        Packet_To_Link_W[21]) );
  FD1LQM1P \Packet_To_Link_W_reg[22]  ( .D(N114), .LD(n68), .CP(Clk_r), .Q(
        Packet_To_Link_W[22]) );
  FD1LQM1P \Packet_To_Link_W_reg[23]  ( .D(N115), .LD(n68), .CP(Clk_r), .Q(
        Packet_To_Link_W[23]) );
  FD1LQM1P \Packet_To_Link_W_reg[26]  ( .D(chosenPacket[26]), .LD(n68), .CP(
        Clk_r), .Q(Packet_To_Link_W[26]) );
  FD1LQM1P \Packet_To_Link_W_reg[28]  ( .D(chosenPacket[28]), .LD(n68), .CP(
        Clk_r), .Q(Packet_To_Link_W[28]) );
  FD1LQM1P \Packet_To_Link_E_reg[31]  ( .D(chosenPacket[31]), .LD(n70), .CP(
        Clk_r), .Q(Packet_To_Link_E[31]) );
  FD1LQM1P \Packet_To_Link_E_reg[30]  ( .D(chosenPacket[30]), .LD(n69), .CP(
        Clk_r), .Q(Packet_To_Link_E[30]) );
  FD1LQM1P \Packet_To_Link_E_reg[29]  ( .D(chosenPacket[29]), .LD(n70), .CP(
        Clk_r), .Q(Packet_To_Link_E[29]) );
  FD1LQM1P \Packet_To_Link_E_reg[27]  ( .D(chosenPacket[27]), .LD(n69), .CP(
        Clk_r), .Q(Packet_To_Link_E[27]) );
  FD1LQM1P \Packet_To_Link_E_reg[25]  ( .D(chosenPacket[25]), .LD(n70), .CP(
        Clk_r), .Q(Packet_To_Link_E[25]) );
  FD1LQM1P \Packet_To_Link_E_reg[16]  ( .D(N108), .LD(n69), .CP(Clk_r), .Q(
        Packet_To_Link_E[16]) );
  FD1LQM1P \Packet_To_Link_E_reg[17]  ( .D(N109), .LD(n70), .CP(Clk_r), .Q(
        Packet_To_Link_E[17]) );
  FD1LQM1P \Packet_To_Link_E_reg[18]  ( .D(N110), .LD(n69), .CP(Clk_r), .Q(
        Packet_To_Link_E[18]) );
  FD1LQM1P \Packet_To_Link_E_reg[19]  ( .D(N111), .LD(n70), .CP(Clk_r), .Q(
        Packet_To_Link_E[19]) );
  FD1LQM1P \Packet_To_Link_E_reg[20]  ( .D(N112), .LD(n69), .CP(Clk_r), .Q(
        Packet_To_Link_E[20]) );
  FD1LQM1P \Packet_To_Link_E_reg[21]  ( .D(N113), .LD(n70), .CP(Clk_r), .Q(
        Packet_To_Link_E[21]) );
  FD1LQM1P \Packet_To_Link_E_reg[22]  ( .D(N114), .LD(n70), .CP(Clk_r), .Q(
        Packet_To_Link_E[22]) );
  FD1LQM1P \Packet_To_Link_E_reg[23]  ( .D(N115), .LD(n70), .CP(Clk_r), .Q(
        Packet_To_Link_E[23]) );
  FD1LQM1P \Packet_To_Link_E_reg[26]  ( .D(chosenPacket[26]), .LD(n70), .CP(
        Clk_r), .Q(Packet_To_Link_E[26]) );
  FD1LQM1P \Packet_To_Link_E_reg[28]  ( .D(chosenPacket[28]), .LD(n70), .CP(
        Clk_r), .Q(Packet_To_Link_E[28]) );
  FD1LQM1P \Packet_To_Link_E_reg[24]  ( .D(chosenPacket[24]), .LD(n70), .CP(
        Clk_r), .Q(Packet_To_Link_E[24]) );
  FD4QM1P \Packet_To_Node_reg[24]  ( .D(n33), .CP(Clk_r), .SD(Rst_n), .Q(
        Packet_To_Node[24]) );
  FD1LQM1P \Packet_To_Link_W_reg[24]  ( .D(chosenPacket[24]), .LD(n68), .CP(
        Clk_r), .Q(Packet_To_Link_W[24]) );
  FD1LQM1P \Packet_To_Link_N_reg[24]  ( .D(chosenPacket[24]), .LD(n39), .CP(
        Clk_r), .Q(Packet_To_Link_N[24]) );
  FD1LQM1P \Packet_To_Link_S_reg[24]  ( .D(chosenPacket[24]), .LD(n40), .CP(
        Clk_r), .Q(Packet_To_Link_S[24]) );
  FD1QM1P \chosenPacket_reg[15]  ( .D(n271), .CP(Clk_r), .Q(chosenPacket[15])
         );
  FD1LQM1P \Packet_To_Link_E_reg[15]  ( .D(chosenPacket[15]), .LD(n70), .CP(
        Clk_r), .Q(Packet_To_Link_E[15]) );
  FD4QM1P \Packet_To_Node_reg[15]  ( .D(n24), .CP(Clk_r), .SD(Rst_n), .Q(
        Packet_To_Node[15]) );
  FD1LQM1P \Packet_To_Link_W_reg[15]  ( .D(chosenPacket[15]), .LD(n68), .CP(
        Clk_r), .Q(Packet_To_Link_W[15]) );
  FD1LQM1P \Packet_To_Link_N_reg[15]  ( .D(chosenPacket[15]), .LD(n39), .CP(
        Clk_r), .Q(Packet_To_Link_N[15]) );
  FD1LQM1P \Packet_To_Link_S_reg[15]  ( .D(chosenPacket[15]), .LD(n40), .CP(
        Clk_r), .Q(Packet_To_Link_S[15]) );
  FD1QM1P \chosenPacket_reg[14]  ( .D(n272), .CP(Clk_r), .Q(chosenPacket[14])
         );
  FD1LQM1P \Packet_To_Link_E_reg[14]  ( .D(chosenPacket[14]), .LD(n70), .CP(
        Clk_r), .Q(Packet_To_Link_E[14]) );
  FD4QM1P \Packet_To_Node_reg[14]  ( .D(n23), .CP(Clk_r), .SD(Rst_n), .Q(
        Packet_To_Node[14]) );
  FD1LQM1P \Packet_To_Link_W_reg[14]  ( .D(chosenPacket[14]), .LD(n68), .CP(
        Clk_r), .Q(Packet_To_Link_W[14]) );
  FD1LQM1P \Packet_To_Link_N_reg[14]  ( .D(chosenPacket[14]), .LD(n39), .CP(
        Clk_r), .Q(Packet_To_Link_N[14]) );
  FD1LQM1P \Packet_To_Link_S_reg[14]  ( .D(chosenPacket[14]), .LD(n40), .CP(
        Clk_r), .Q(Packet_To_Link_S[14]) );
  FD1QM1P \chosenPacket_reg[13]  ( .D(n273), .CP(Clk_r), .Q(chosenPacket[13])
         );
  FD1LQM1P \Packet_To_Link_E_reg[13]  ( .D(chosenPacket[13]), .LD(n70), .CP(
        Clk_r), .Q(Packet_To_Link_E[13]) );
  FD4QM1P \Packet_To_Node_reg[13]  ( .D(n22), .CP(Clk_r), .SD(Rst_n), .Q(
        Packet_To_Node[13]) );
  FD1LQM1P \Packet_To_Link_W_reg[13]  ( .D(chosenPacket[13]), .LD(n68), .CP(
        Clk_r), .Q(Packet_To_Link_W[13]) );
  FD1LQM1P \Packet_To_Link_N_reg[13]  ( .D(chosenPacket[13]), .LD(n39), .CP(
        Clk_r), .Q(Packet_To_Link_N[13]) );
  FD1LQM1P \Packet_To_Link_S_reg[13]  ( .D(chosenPacket[13]), .LD(n40), .CP(
        Clk_r), .Q(Packet_To_Link_S[13]) );
  FD1QM1P \chosenPacket_reg[12]  ( .D(n274), .CP(Clk_r), .Q(chosenPacket[12])
         );
  FD1LQM1P \Packet_To_Link_E_reg[12]  ( .D(chosenPacket[12]), .LD(n70), .CP(
        Clk_r), .Q(Packet_To_Link_E[12]) );
  FD4QM1P \Packet_To_Node_reg[12]  ( .D(n21), .CP(Clk_r), .SD(Rst_n), .Q(
        Packet_To_Node[12]) );
  FD1LQM1P \Packet_To_Link_W_reg[12]  ( .D(chosenPacket[12]), .LD(n68), .CP(
        Clk_r), .Q(Packet_To_Link_W[12]) );
  FD1LQM1P \Packet_To_Link_N_reg[12]  ( .D(chosenPacket[12]), .LD(n39), .CP(
        Clk_r), .Q(Packet_To_Link_N[12]) );
  FD1LQM1P \Packet_To_Link_S_reg[12]  ( .D(chosenPacket[12]), .LD(n40), .CP(
        Clk_r), .Q(Packet_To_Link_S[12]) );
  FD1QM1P \chosenPacket_reg[11]  ( .D(n275), .CP(Clk_r), .Q(chosenPacket[11])
         );
  FD1LQM1P \Packet_To_Link_E_reg[11]  ( .D(chosenPacket[11]), .LD(n70), .CP(
        Clk_r), .Q(Packet_To_Link_E[11]) );
  FD4QM1P \Packet_To_Node_reg[11]  ( .D(n20), .CP(Clk_r), .SD(Rst_n), .Q(
        Packet_To_Node[11]) );
  FD1LQM1P \Packet_To_Link_W_reg[11]  ( .D(chosenPacket[11]), .LD(n68), .CP(
        Clk_r), .Q(Packet_To_Link_W[11]) );
  FD1LQM1P \Packet_To_Link_N_reg[11]  ( .D(chosenPacket[11]), .LD(n39), .CP(
        Clk_r), .Q(Packet_To_Link_N[11]) );
  FD1LQM1P \Packet_To_Link_S_reg[11]  ( .D(chosenPacket[11]), .LD(n40), .CP(
        Clk_r), .Q(Packet_To_Link_S[11]) );
  FD1QM1P \chosenPacket_reg[10]  ( .D(n276), .CP(Clk_r), .Q(chosenPacket[10])
         );
  FD1LQM1P \Packet_To_Link_E_reg[10]  ( .D(chosenPacket[10]), .LD(n69), .CP(
        Clk_r), .Q(Packet_To_Link_E[10]) );
  FD4QM1P \Packet_To_Node_reg[10]  ( .D(n19), .CP(Clk_r), .SD(Rst_n), .Q(
        Packet_To_Node[10]) );
  FD1LQM1P \Packet_To_Link_W_reg[10]  ( .D(chosenPacket[10]), .LD(n67), .CP(
        Clk_r), .Q(Packet_To_Link_W[10]) );
  FD1LQM1P \Packet_To_Link_N_reg[10]  ( .D(chosenPacket[10]), .LD(n39), .CP(
        Clk_r), .Q(Packet_To_Link_N[10]) );
  FD1LQM1P \Packet_To_Link_S_reg[10]  ( .D(chosenPacket[10]), .LD(n40), .CP(
        Clk_r), .Q(Packet_To_Link_S[10]) );
  FD1QM1P \chosenPacket_reg[9]  ( .D(n277), .CP(Clk_r), .Q(chosenPacket[9]) );
  FD1LQM1P \Packet_To_Link_E_reg[9]  ( .D(chosenPacket[9]), .LD(n69), .CP(
        Clk_r), .Q(Packet_To_Link_E[9]) );
  FD4QM1P \Packet_To_Node_reg[9]  ( .D(n18), .CP(Clk_r), .SD(Rst_n), .Q(
        Packet_To_Node[9]) );
  FD1LQM1P \Packet_To_Link_W_reg[9]  ( .D(chosenPacket[9]), .LD(n67), .CP(
        Clk_r), .Q(Packet_To_Link_W[9]) );
  FD1LQM1P \Packet_To_Link_N_reg[9]  ( .D(chosenPacket[9]), .LD(n39), .CP(
        Clk_r), .Q(Packet_To_Link_N[9]) );
  FD1LQM1P \Packet_To_Link_S_reg[9]  ( .D(chosenPacket[9]), .LD(n40), .CP(
        Clk_r), .Q(Packet_To_Link_S[9]) );
  FD1QM1P \chosenPacket_reg[8]  ( .D(n278), .CP(Clk_r), .Q(chosenPacket[8]) );
  FD1LQM1P \Packet_To_Link_E_reg[8]  ( .D(chosenPacket[8]), .LD(n69), .CP(
        Clk_r), .Q(Packet_To_Link_E[8]) );
  FD4QM1P \Packet_To_Node_reg[8]  ( .D(n17), .CP(Clk_r), .SD(Rst_n), .Q(
        Packet_To_Node[8]) );
  FD1LQM1P \Packet_To_Link_W_reg[8]  ( .D(chosenPacket[8]), .LD(n67), .CP(
        Clk_r), .Q(Packet_To_Link_W[8]) );
  FD1LQM1P \Packet_To_Link_N_reg[8]  ( .D(chosenPacket[8]), .LD(n39), .CP(
        Clk_r), .Q(Packet_To_Link_N[8]) );
  FD1LQM1P \Packet_To_Link_S_reg[8]  ( .D(chosenPacket[8]), .LD(n40), .CP(
        Clk_r), .Q(Packet_To_Link_S[8]) );
  FD1QM1P \chosenPacket_reg[7]  ( .D(n279), .CP(Clk_r), .Q(chosenPacket[7]) );
  FD1LQM1P \Packet_To_Link_E_reg[7]  ( .D(chosenPacket[7]), .LD(n69), .CP(
        Clk_r), .Q(Packet_To_Link_E[7]) );
  FD4QM1P \Packet_To_Node_reg[7]  ( .D(n16), .CP(Clk_r), .SD(Rst_n), .Q(
        Packet_To_Node[7]) );
  FD1LQM1P \Packet_To_Link_W_reg[7]  ( .D(chosenPacket[7]), .LD(n67), .CP(
        Clk_r), .Q(Packet_To_Link_W[7]) );
  FD1LQM1P \Packet_To_Link_N_reg[7]  ( .D(chosenPacket[7]), .LD(n39), .CP(
        Clk_r), .Q(Packet_To_Link_N[7]) );
  FD1LQM1P \Packet_To_Link_S_reg[7]  ( .D(chosenPacket[7]), .LD(n40), .CP(
        Clk_r), .Q(Packet_To_Link_S[7]) );
  FD1QM1P \chosenPacket_reg[6]  ( .D(n280), .CP(Clk_r), .Q(chosenPacket[6]) );
  FD1LQM1P \Packet_To_Link_E_reg[6]  ( .D(chosenPacket[6]), .LD(n69), .CP(
        Clk_r), .Q(Packet_To_Link_E[6]) );
  FD4QM1P \Packet_To_Node_reg[6]  ( .D(n15), .CP(Clk_r), .SD(Rst_n), .Q(
        Packet_To_Node[6]) );
  FD1LQM1P \Packet_To_Link_W_reg[6]  ( .D(chosenPacket[6]), .LD(n67), .CP(
        Clk_r), .Q(Packet_To_Link_W[6]) );
  FD1LQM1P \Packet_To_Link_N_reg[6]  ( .D(chosenPacket[6]), .LD(n39), .CP(
        Clk_r), .Q(Packet_To_Link_N[6]) );
  FD1LQM1P \Packet_To_Link_S_reg[6]  ( .D(chosenPacket[6]), .LD(n40), .CP(
        Clk_r), .Q(Packet_To_Link_S[6]) );
  FD1QM1P \chosenPacket_reg[5]  ( .D(n281), .CP(Clk_r), .Q(chosenPacket[5]) );
  FD1LQM1P \Packet_To_Link_E_reg[5]  ( .D(chosenPacket[5]), .LD(n69), .CP(
        Clk_r), .Q(Packet_To_Link_E[5]) );
  FD4QM1P \Packet_To_Node_reg[5]  ( .D(n14), .CP(Clk_r), .SD(Rst_n), .Q(
        Packet_To_Node[5]) );
  FD1LQM1P \Packet_To_Link_W_reg[5]  ( .D(chosenPacket[5]), .LD(n67), .CP(
        Clk_r), .Q(Packet_To_Link_W[5]) );
  FD1LQM1P \Packet_To_Link_N_reg[5]  ( .D(chosenPacket[5]), .LD(n39), .CP(
        Clk_r), .Q(Packet_To_Link_N[5]) );
  FD1LQM1P \Packet_To_Link_S_reg[5]  ( .D(chosenPacket[5]), .LD(n40), .CP(
        Clk_r), .Q(Packet_To_Link_S[5]) );
  FD1QM1P \chosenPacket_reg[4]  ( .D(n282), .CP(Clk_r), .Q(chosenPacket[4]) );
  FD1LQM1P \Packet_To_Link_E_reg[4]  ( .D(chosenPacket[4]), .LD(n69), .CP(
        Clk_r), .Q(Packet_To_Link_E[4]) );
  FD4QM1P \Packet_To_Node_reg[4]  ( .D(n13), .CP(Clk_r), .SD(Rst_n), .Q(
        Packet_To_Node[4]) );
  FD1LQM1P \Packet_To_Link_W_reg[4]  ( .D(chosenPacket[4]), .LD(n67), .CP(
        Clk_r), .Q(Packet_To_Link_W[4]) );
  FD1LQM1P \Packet_To_Link_N_reg[4]  ( .D(chosenPacket[4]), .LD(n39), .CP(
        Clk_r), .Q(Packet_To_Link_N[4]) );
  FD1LQM1P \Packet_To_Link_S_reg[4]  ( .D(chosenPacket[4]), .LD(n40), .CP(
        Clk_r), .Q(Packet_To_Link_S[4]) );
  FD1QM1P \chosenPacket_reg[3]  ( .D(n283), .CP(Clk_r), .Q(chosenPacket[3]) );
  FD1LQM1P \Packet_To_Link_E_reg[3]  ( .D(chosenPacket[3]), .LD(n69), .CP(
        Clk_r), .Q(Packet_To_Link_E[3]) );
  FD4QM1P \Packet_To_Node_reg[3]  ( .D(n12), .CP(Clk_r), .SD(Rst_n), .Q(
        Packet_To_Node[3]) );
  FD1LQM1P \Packet_To_Link_W_reg[3]  ( .D(chosenPacket[3]), .LD(n67), .CP(
        Clk_r), .Q(Packet_To_Link_W[3]) );
  FD1LQM1P \Packet_To_Link_N_reg[3]  ( .D(chosenPacket[3]), .LD(n39), .CP(
        Clk_r), .Q(Packet_To_Link_N[3]) );
  FD1LQM1P \Packet_To_Link_S_reg[3]  ( .D(chosenPacket[3]), .LD(n40), .CP(
        Clk_r), .Q(Packet_To_Link_S[3]) );
  FD1QM1P \chosenPacket_reg[2]  ( .D(n284), .CP(Clk_r), .Q(chosenPacket[2]) );
  FD1LQM1P \Packet_To_Link_E_reg[2]  ( .D(chosenPacket[2]), .LD(n69), .CP(
        Clk_r), .Q(Packet_To_Link_E[2]) );
  FD4QM1P \Packet_To_Node_reg[2]  ( .D(n11), .CP(Clk_r), .SD(Rst_n), .Q(
        Packet_To_Node[2]) );
  FD1LQM1P \Packet_To_Link_W_reg[2]  ( .D(chosenPacket[2]), .LD(n67), .CP(
        Clk_r), .Q(Packet_To_Link_W[2]) );
  FD1LQM1P \Packet_To_Link_N_reg[2]  ( .D(chosenPacket[2]), .LD(n39), .CP(
        Clk_r), .Q(Packet_To_Link_N[2]) );
  FD1LQM1P \Packet_To_Link_S_reg[2]  ( .D(chosenPacket[2]), .LD(n40), .CP(
        Clk_r), .Q(Packet_To_Link_S[2]) );
  FD1QM1P \chosenPacket_reg[1]  ( .D(n285), .CP(Clk_r), .Q(chosenPacket[1]) );
  FD1LQM1P \Packet_To_Link_E_reg[1]  ( .D(chosenPacket[1]), .LD(n69), .CP(
        Clk_r), .Q(Packet_To_Link_E[1]) );
  FD4QM1P \Packet_To_Node_reg[1]  ( .D(n10), .CP(Clk_r), .SD(Rst_n), .Q(
        Packet_To_Node[1]) );
  FD1LQM1P \Packet_To_Link_W_reg[1]  ( .D(chosenPacket[1]), .LD(n67), .CP(
        Clk_r), .Q(Packet_To_Link_W[1]) );
  FD1LQM1P \Packet_To_Link_N_reg[1]  ( .D(chosenPacket[1]), .LD(n39), .CP(
        Clk_r), .Q(Packet_To_Link_N[1]) );
  FD1LQM1P \Packet_To_Link_S_reg[1]  ( .D(chosenPacket[1]), .LD(n40), .CP(
        Clk_r), .Q(Packet_To_Link_S[1]) );
  FD1QM1P \chosenPacket_reg[0]  ( .D(n286), .CP(Clk_r), .Q(chosenPacket[0]) );
  FD1LQM1P \Packet_To_Link_E_reg[0]  ( .D(chosenPacket[0]), .LD(n69), .CP(
        Clk_r), .Q(Packet_To_Link_E[0]) );
  FD4QM1P \Packet_To_Node_reg[0]  ( .D(n9), .CP(Clk_r), .SD(Rst_n), .Q(
        Packet_To_Node[0]) );
  FD1LQM1P \Packet_To_Link_W_reg[0]  ( .D(chosenPacket[0]), .LD(n67), .CP(
        Clk_r), .Q(Packet_To_Link_W[0]) );
  FD1LQM1P \Packet_To_Link_N_reg[0]  ( .D(chosenPacket[0]), .LD(n39), .CP(
        Clk_r), .Q(Packet_To_Link_N[0]) );
  FD1LQM1P \Packet_To_Link_S_reg[0]  ( .D(chosenPacket[0]), .LD(n40), .CP(
        Clk_r), .Q(Packet_To_Link_S[0]) );
  FD1QM1P \chosenPacket_reg[23]  ( .D(n262), .CP(Clk_r), .Q(chosenPacket[23])
         );
  FD1QM1P \chosenPacket_reg[16]  ( .D(n260), .CP(Clk_r), .Q(chosenPacket[16])
         );
  FD1QM1P \chosenPacket_reg[17]  ( .D(n259), .CP(Clk_r), .Q(chosenPacket[17])
         );
  FD1QM1P \chosenPacket_reg[18]  ( .D(n258), .CP(Clk_r), .Q(chosenPacket[18])
         );
  FD1QM1P \chosenPacket_reg[19]  ( .D(n257), .CP(Clk_r), .Q(chosenPacket[19])
         );
  FD1QM1P \chosenPacket_reg[20]  ( .D(n256), .CP(Clk_r), .Q(chosenPacket[20])
         );
  FD1QM1P \chosenPacket_reg[21]  ( .D(n255), .CP(Clk_r), .Q(chosenPacket[21])
         );
  FD1QM1P \chosenPacket_reg[22]  ( .D(n254), .CP(Clk_r), .Q(chosenPacket[22])
         );
  FD4QM1P \TxQueue_Write_reg[0]  ( .D(n53), .CP(Clk_r), .SD(Rst_n), .Q(n54) );
  FD4QM1P \RxQueue_Read_reg[1]  ( .D(n226), .CP(Clk_r), .SD(Rst_n), .Q(n52) );
  FD4QM1P \nextStage_reg[0]  ( .D(n7), .CP(Clk_r), .SD(Rst_n), .Q(n8) );
  FD2QM1P \TxQueue_Write_reg[3]  ( .D(n253), .CP(Clk_r), .CD(Rst_n), .Q(
        TxQueue_Write_N) );
  FD2QM1P \TxQueue_Write_reg[2]  ( .D(n252), .CP(Clk_r), .CD(Rst_n), .Q(
        TxQueue_Write_S) );
  FD2QM1P To_Node_Write_reg ( .D(n261), .CP(Clk_r), .CD(Rst_n), .Q(
        To_Node_Write) );
  FD2QM1P \TxQueue_Write_reg[1]  ( .D(n251), .CP(Clk_r), .CD(Rst_n), .Q(
        TxQueue_Write_W) );
  FD2QM1P \RxQueue_Read_reg[2]  ( .D(n247), .CP(Clk_r), .CD(Rst_n), .Q(
        RxQueue_Read_S) );
  FD2QM1P \RxQueue_Read_reg[0]  ( .D(n249), .CP(Clk_r), .CD(Rst_n), .Q(
        RxQueue_Read_E) );
  FD2QM1P \RxQueue_Read_reg[3]  ( .D(n246), .CP(Clk_r), .CD(Rst_n), .Q(
        RxQueue_Read_N) );
  FD2QM1P \RxQueue_Read_reg[4]  ( .D(n245), .CP(Clk_r), .CD(Rst_n), .Q(
        Node_Read) );
  FD2LQM1P \Packet_To_Node_reg[22]  ( .D(n48), .LD(n107), .CP(Clk_r), .CD(
        Rst_n), .Q(n49) );
  BUFM2P U3 ( .A(n192), .Z(n64) );
  BUFM2P U4 ( .A(n192), .Z(n63) );
  BUFM2P U5 ( .A(n156), .Z(n51) );
  ND2M2P U6 ( .A(n305), .B(Rst_n), .Z(n155) );
  AND2M1P U7 ( .A(n223), .B(Rst_n), .Z(n233) );
  NR2M1P U8 ( .A(n227), .B(n155), .Z(n191) );
  AOI211M1P U9 ( .A(n43), .B(Router_Address[5]), .C(Router_Address[4]), .D(
        n236), .Z(n31) );
  N1M1P U10 ( .A(n222), .Z(n36) );
  OAI22CDNM1P U11 ( .A(n31), .B(n36), .C(Router_Address[6]), .D(n42), .Z(n46)
         );
  MAJN3M1P U12 ( .A(n41), .B(Router_Address[7]), .C(n46), .Z(n47) );
  ND3CNM1P U13 ( .C(TxQueue_Full_E), .A(Link_Config[0]), .B(n47), .Z(n302) );
  NR2FM2P U14 ( .A(n228), .B(n155), .Z(n189) );
  NR2FM3P U15 ( .A(n57), .B(n155), .Z(n156) );
  BUFM8P U16 ( .A(n189), .Z(n56) );
  N1M2P U17 ( .A(n107), .Z(n66) );
  NR2BNM2P U18 ( .B(n307), .A(To_Node_Full), .Z(n107) );
  N1M1P U19 ( .A(n49), .Z(Packet_To_Node[22]) );
  N1M1P U20 ( .A(N114), .Z(n48) );
  BUFM3P U21 ( .A(n190), .Z(n50) );
  NR2M1P U22 ( .A(dataLocation[0]), .B(n80), .Z(N43) );
  N1M1P U23 ( .A(n54), .Z(TxQueue_Write_E) );
  N1M2P U24 ( .A(n52), .Z(RxQueue_Read_W) );
  N1M1P U25 ( .A(n8), .Z(n223) );
  N1M1P U26 ( .A(n6), .Z(n80) );
  N1M2P U27 ( .A(n66), .Z(n65) );
  AND2M4P U28 ( .A(n233), .B(n231), .Z(n39) );
  AND2M4P U29 ( .A(n230), .B(n233), .Z(n40) );
  BUFM2P U30 ( .A(n155), .Z(n55) );
  MUX21LM1P U31 ( .A(chosenPacket[23]), .B(n79), .S(n78), .Z(N115) );
  N1M1P U32 ( .A(chosenPacket[31]), .Z(n41) );
  MUX21LM1P U33 ( .A(chosenPacket[22]), .B(n71), .S(n77), .Z(N114) );
  BUFM2P U34 ( .A(n37), .Z(n70) );
  BUFM2P U35 ( .A(n37), .Z(n69) );
  BUFM2P U36 ( .A(n38), .Z(n68) );
  BUFM2P U37 ( .A(n38), .Z(n67) );
  BUFM2P U38 ( .A(n191), .Z(n59) );
  BUFM2P U39 ( .A(n191), .Z(n60) );
  BUFM2P U40 ( .A(n191), .Z(n61) );
  BUFM2P U41 ( .A(n190), .Z(n58) );
  NR2FM1P U42 ( .A(n223), .B(n160), .Z(n305) );
  N1M1P U43 ( .A(n250), .Z(n53) );
  BUFM1P U44 ( .A(n191), .Z(n62) );
  NR2BNM1P U45 ( .B(n225), .A(n155), .Z(n190) );
  ND3M1P U46 ( .A(n84), .B(n83), .C(n82), .Z(n160) );
  AOI22DNM1P U47 ( .A(n81), .B(RxQueue_Empty_S), .D(n57), .C(Node_Queue_Empty), 
        .Z(n83) );
  MUX41HM3P U48 ( .D0(Link_Config[0]), .D1(Link_Config[2]), .D2(Link_Config[1]), .D3(Link_Config[3]), .A(N44), .B(N43), .Z(N48) );
  NR2M1P U49 ( .A(n6), .B(n155), .Z(n192) );
  AOI22DNM1P U50 ( .A(n225), .B(RxQueue_Empty_W), .D(n228), .C(RxQueue_Empty_N), .Z(n82) );
  N1M1P U51 ( .A(chosenPacket[22]), .Z(n71) );
  N1M1P U52 ( .A(chosenPacket[20]), .Z(n73) );
  AND3M1P U53 ( .A(chosenPacket[16]), .B(chosenPacket[17]), .C(
        chosenPacket[18]), .Z(n76) );
  ND2M1P U54 ( .A(n76), .B(chosenPacket[19]), .Z(n74) );
  NR2M1P U55 ( .A(n73), .B(n74), .Z(n72) );
  ND2M1P U56 ( .A(n72), .B(chosenPacket[21]), .Z(n77) );
  OR2M1P U57 ( .A(n72), .B(chosenPacket[21]), .Z(n196) );
  ND2M1P U58 ( .A(n77), .B(n196), .Z(n240) );
  N1M1P U59 ( .A(n240), .Z(N113) );
  AOI21M1P U60 ( .A(n74), .B(n73), .C(n72), .Z(N112) );
  OAI21M1P U61 ( .A(n76), .B(chosenPacket[19]), .C(n74), .Z(n242) );
  N1M1P U62 ( .A(n242), .Z(N111) );
  AOI21M1P U63 ( .A(chosenPacket[17]), .B(chosenPacket[16]), .C(
        chosenPacket[18]), .Z(n75) );
  NR2M1P U64 ( .A(n76), .B(n75), .Z(N110) );
  OAI22CDNM1P U65 ( .A(chosenPacket[17]), .B(chosenPacket[16]), .C(
        chosenPacket[16]), .D(chosenPacket[17]), .Z(n244) );
  N1M1P U66 ( .A(n244), .Z(N109) );
  N1M1P U67 ( .A(chosenPacket[16]), .Z(N108) );
  N1M1P U68 ( .A(chosenPacket[23]), .Z(n79) );
  ND2BNM1P U69 ( .B(n77), .A(chosenPacket[22]), .Z(n78) );
  N1M1P U70 ( .A(chosenPacket[25]), .Z(n45) );
  N1M1P U71 ( .A(chosenPacket[27]), .Z(n44) );
  N1M1P U72 ( .A(chosenPacket[29]), .Z(n43) );
  N1M1P U73 ( .A(chosenPacket[30]), .Z(n42) );
  ND3M1P U74 ( .A(dataLocation[0]), .B(n6), .C(dataLocation[1]), .Z(n57) );
  ND2M1P U75 ( .A(N43), .B(dataLocation[1]), .Z(n228) );
  NR3CNM1P U76 ( .C(dataLocation[0]), .A(dataLocation[1]), .B(n80), .Z(n81) );
  N1M1P U77 ( .A(n81), .Z(n227) );
  ND2M1P U78 ( .A(n228), .B(n227), .Z(N44) );
  AOI22DNM1P U79 ( .A(RxQueue_Empty_E), .B(n80), .D(N48), .C(n57), .Z(n84) );
  NR2BNM1P U80 ( .B(N43), .A(dataLocation[1]), .Z(n225) );
  AOI22M1P U81 ( .A(Packet_From_Link_E[0]), .B(n64), .C(chosenPacket[0]), .D(
        n55), .Z(n87) );
  AOI22M1P U82 ( .A(n189), .B(Packet_From_Link_N[0]), .C(n59), .D(
        Packet_From_Link_S[0]), .Z(n86) );
  AOI22M1P U83 ( .A(n50), .B(Packet_From_Link_W[0]), .C(n156), .D(
        Packet_From_Node[0]), .Z(n85) );
  ND3M1P U84 ( .A(n87), .B(n86), .C(n85), .Z(n286) );
  AOI22M1P U85 ( .A(Packet_From_Link_E[1]), .B(n63), .C(chosenPacket[1]), .D(
        n55), .Z(n90) );
  AOI22M1P U86 ( .A(n189), .B(Packet_From_Link_N[1]), .C(n59), .D(
        Packet_From_Link_S[1]), .Z(n89) );
  AOI22M1P U87 ( .A(n58), .B(Packet_From_Link_W[1]), .C(n156), .D(
        Packet_From_Node[1]), .Z(n88) );
  ND3M1P U88 ( .A(n90), .B(n89), .C(n88), .Z(n285) );
  AOI22M1P U89 ( .A(Packet_From_Link_E[2]), .B(n63), .C(chosenPacket[2]), .D(
        n55), .Z(n93) );
  AOI22M1P U90 ( .A(n189), .B(Packet_From_Link_N[2]), .C(n59), .D(
        Packet_From_Link_S[2]), .Z(n92) );
  AOI22M1P U91 ( .A(n50), .B(Packet_From_Link_W[2]), .C(n156), .D(
        Packet_From_Node[2]), .Z(n91) );
  ND3M1P U92 ( .A(n93), .B(n92), .C(n91), .Z(n284) );
  AOI22M1P U93 ( .A(Packet_From_Link_E[3]), .B(n64), .C(chosenPacket[3]), .D(
        n55), .Z(n96) );
  AOI22M1P U94 ( .A(n189), .B(Packet_From_Link_N[3]), .C(n59), .D(
        Packet_From_Link_S[3]), .Z(n95) );
  AOI22M1P U95 ( .A(n50), .B(Packet_From_Link_W[3]), .C(n156), .D(
        Packet_From_Node[3]), .Z(n94) );
  ND3M1P U96 ( .A(n96), .B(n95), .C(n94), .Z(n283) );
  AOI22M1P U97 ( .A(Packet_From_Link_E[4]), .B(n63), .C(chosenPacket[4]), .D(
        n55), .Z(n99) );
  AOI22M1P U98 ( .A(n189), .B(Packet_From_Link_N[4]), .C(n59), .D(
        Packet_From_Link_S[4]), .Z(n98) );
  AOI22M1P U99 ( .A(n50), .B(Packet_From_Link_W[4]), .C(n156), .D(
        Packet_From_Node[4]), .Z(n97) );
  ND3M1P U100 ( .A(n99), .B(n98), .C(n97), .Z(n282) );
  AOI22M1P U101 ( .A(Packet_From_Link_E[5]), .B(n64), .C(chosenPacket[5]), .D(
        n55), .Z(n102) );
  AOI22M1P U102 ( .A(n189), .B(Packet_From_Link_N[5]), .C(n59), .D(
        Packet_From_Link_S[5]), .Z(n101) );
  AOI22M1P U103 ( .A(n50), .B(Packet_From_Link_W[5]), .C(n51), .D(
        Packet_From_Node[5]), .Z(n100) );
  ND3M1P U104 ( .A(n102), .B(n101), .C(n100), .Z(n281) );
  AOI22M1P U105 ( .A(Packet_From_Link_E[6]), .B(n63), .C(chosenPacket[6]), .D(
        n55), .Z(n105) );
  AOI22M1P U106 ( .A(n189), .B(Packet_From_Link_N[6]), .C(n59), .D(
        Packet_From_Link_S[6]), .Z(n104) );
  AOI22M1P U107 ( .A(n50), .B(Packet_From_Link_W[6]), .C(n51), .D(
        Packet_From_Node[6]), .Z(n103) );
  ND3M1P U108 ( .A(n105), .B(n104), .C(n103), .Z(n280) );
  AOI22M1P U109 ( .A(Packet_From_Link_E[7]), .B(n64), .C(chosenPacket[7]), .D(
        n55), .Z(n109) );
  AOI22M1P U110 ( .A(n189), .B(Packet_From_Link_N[7]), .C(n59), .D(
        Packet_From_Link_S[7]), .Z(n108) );
  AOI22M1P U111 ( .A(n50), .B(Packet_From_Link_W[7]), .C(n51), .D(
        Packet_From_Node[7]), .Z(n106) );
  ND3M1P U112 ( .A(n109), .B(n108), .C(n106), .Z(n279) );
  AOI22M1P U113 ( .A(Packet_From_Link_E[8]), .B(n63), .C(chosenPacket[8]), .D(
        n55), .Z(n112) );
  AOI22M1P U114 ( .A(n189), .B(Packet_From_Link_N[8]), .C(n59), .D(
        Packet_From_Link_S[8]), .Z(n111) );
  AOI22M1P U115 ( .A(n50), .B(Packet_From_Link_W[8]), .C(n51), .D(
        Packet_From_Node[8]), .Z(n110) );
  ND3M1P U116 ( .A(n112), .B(n111), .C(n110), .Z(n278) );
  AOI22M1P U117 ( .A(Packet_From_Link_E[9]), .B(n64), .C(chosenPacket[9]), .D(
        n55), .Z(n115) );
  AOI22M1P U118 ( .A(n56), .B(Packet_From_Link_N[9]), .C(n59), .D(
        Packet_From_Link_S[9]), .Z(n114) );
  AOI22M1P U119 ( .A(n50), .B(Packet_From_Link_W[9]), .C(n51), .D(
        Packet_From_Node[9]), .Z(n113) );
  ND3M1P U120 ( .A(n115), .B(n114), .C(n113), .Z(n277) );
  AOI22M1P U121 ( .A(Packet_From_Link_E[10]), .B(n63), .C(chosenPacket[10]), 
        .D(n55), .Z(n118) );
  AOI22M1P U122 ( .A(n56), .B(Packet_From_Link_N[10]), .C(n60), .D(
        Packet_From_Link_S[10]), .Z(n117) );
  AOI22M1P U123 ( .A(n50), .B(Packet_From_Link_W[10]), .C(n51), .D(
        Packet_From_Node[10]), .Z(n116) );
  ND3M1P U124 ( .A(n118), .B(n117), .C(n116), .Z(n276) );
  AOI22M1P U125 ( .A(Packet_From_Link_E[11]), .B(n64), .C(chosenPacket[11]), 
        .D(n55), .Z(n121) );
  AOI22M1P U126 ( .A(n56), .B(Packet_From_Link_N[11]), .C(n60), .D(
        Packet_From_Link_S[11]), .Z(n120) );
  AOI22M1P U127 ( .A(n50), .B(Packet_From_Link_W[11]), .C(n51), .D(
        Packet_From_Node[11]), .Z(n119) );
  ND3M1P U128 ( .A(n121), .B(n120), .C(n119), .Z(n275) );
  AOI22M1P U129 ( .A(Packet_From_Link_E[12]), .B(n64), .C(chosenPacket[12]), 
        .D(n55), .Z(n124) );
  AOI22M1P U130 ( .A(n56), .B(Packet_From_Link_N[12]), .C(n60), .D(
        Packet_From_Link_S[12]), .Z(n123) );
  AOI22M1P U131 ( .A(n50), .B(Packet_From_Link_W[12]), .C(n51), .D(
        Packet_From_Node[12]), .Z(n122) );
  ND3M1P U132 ( .A(n124), .B(n123), .C(n122), .Z(n274) );
  AOI22M1P U133 ( .A(Packet_From_Link_E[13]), .B(n64), .C(chosenPacket[13]), 
        .D(n55), .Z(n127) );
  AOI22M1P U134 ( .A(n56), .B(Packet_From_Link_N[13]), .C(n60), .D(
        Packet_From_Link_S[13]), .Z(n126) );
  AOI22M1P U135 ( .A(n50), .B(Packet_From_Link_W[13]), .C(n51), .D(
        Packet_From_Node[13]), .Z(n125) );
  ND3M1P U136 ( .A(n127), .B(n126), .C(n125), .Z(n273) );
  AOI22M1P U137 ( .A(Packet_From_Link_E[14]), .B(n64), .C(chosenPacket[14]), 
        .D(n55), .Z(n130) );
  AOI22M1P U138 ( .A(n56), .B(Packet_From_Link_N[14]), .C(n60), .D(
        Packet_From_Link_S[14]), .Z(n129) );
  AOI22M1P U139 ( .A(n50), .B(Packet_From_Link_W[14]), .C(n51), .D(
        Packet_From_Node[14]), .Z(n128) );
  ND3M1P U140 ( .A(n130), .B(n129), .C(n128), .Z(n272) );
  AOI22M1P U141 ( .A(Packet_From_Link_E[15]), .B(n64), .C(chosenPacket[15]), 
        .D(n55), .Z(n133) );
  AOI22M1P U142 ( .A(n56), .B(Packet_From_Link_N[15]), .C(n60), .D(
        Packet_From_Link_S[15]), .Z(n132) );
  AOI22M1P U143 ( .A(n50), .B(Packet_From_Link_W[15]), .C(n51), .D(
        Packet_From_Node[15]), .Z(n131) );
  ND3M1P U144 ( .A(n133), .B(n132), .C(n131), .Z(n271) );
  AOI22M1P U145 ( .A(chosenPacket[24]), .B(n55), .C(n64), .D(
        Packet_From_Link_E[24]), .Z(n136) );
  AOI22M1P U146 ( .A(n56), .B(Packet_From_Link_N[24]), .C(n60), .D(
        Packet_From_Link_S[24]), .Z(n135) );
  AOI22M1P U147 ( .A(n50), .B(Packet_From_Link_W[24]), .C(n51), .D(
        Packet_From_Node_24), .Z(n134) );
  ND3M1P U148 ( .A(n136), .B(n135), .C(n134), .Z(n270) );
  AOI22M1P U149 ( .A(chosenPacket[25]), .B(n55), .C(n64), .D(
        Packet_From_Link_E[25]), .Z(n139) );
  AOI22M1P U150 ( .A(n56), .B(Packet_From_Link_N[25]), .C(n60), .D(
        Packet_From_Link_S[25]), .Z(n138) );
  AOI22M1P U151 ( .A(n50), .B(Packet_From_Link_W[25]), .C(n51), .D(
        Packet_From_Node_25), .Z(n137) );
  ND3M1P U152 ( .A(n139), .B(n138), .C(n137), .Z(n269) );
  AOI22M1P U153 ( .A(chosenPacket[26]), .B(n55), .C(n64), .D(
        Packet_From_Link_E[26]), .Z(n142) );
  AOI22M1P U154 ( .A(n56), .B(Packet_From_Link_N[26]), .C(n60), .D(
        Packet_From_Link_S[26]), .Z(n141) );
  AOI22M1P U155 ( .A(n50), .B(Packet_From_Link_W[26]), .C(n51), .D(
        Packet_From_Node_26), .Z(n140) );
  ND3M1P U156 ( .A(n142), .B(n141), .C(n140), .Z(n268) );
  AOI22M1P U157 ( .A(chosenPacket[27]), .B(n55), .C(n64), .D(
        Packet_From_Link_E[27]), .Z(n145) );
  AOI22M1P U158 ( .A(n56), .B(Packet_From_Link_N[27]), .C(n60), .D(
        Packet_From_Link_S[27]), .Z(n144) );
  AOI22M1P U159 ( .A(n50), .B(Packet_From_Link_W[27]), .C(n51), .D(
        Packet_From_Node_27), .Z(n143) );
  ND3M1P U160 ( .A(n145), .B(n144), .C(n143), .Z(n267) );
  AOI22M1P U161 ( .A(chosenPacket[28]), .B(n55), .C(n64), .D(
        Packet_From_Link_E[28]), .Z(n148) );
  AOI22M1P U162 ( .A(n56), .B(Packet_From_Link_N[28]), .C(n61), .D(
        Packet_From_Link_S[28]), .Z(n147) );
  AOI22M1P U163 ( .A(n58), .B(Packet_From_Link_W[28]), .C(n51), .D(
        Packet_From_Node_28), .Z(n146) );
  ND3M1P U164 ( .A(n148), .B(n147), .C(n146), .Z(n266) );
  AOI22M1P U165 ( .A(chosenPacket[29]), .B(n55), .C(n64), .D(
        Packet_From_Link_E[29]), .Z(n151) );
  AOI22M1P U166 ( .A(n56), .B(Packet_From_Link_N[29]), .C(n61), .D(
        Packet_From_Link_S[29]), .Z(n150) );
  AOI22M1P U167 ( .A(n58), .B(Packet_From_Link_W[29]), .C(n51), .D(
        Packet_From_Node_29), .Z(n149) );
  ND3M1P U168 ( .A(n151), .B(n150), .C(n149), .Z(n265) );
  AOI22M1P U169 ( .A(chosenPacket[30]), .B(n55), .C(n63), .D(
        Packet_From_Link_E[30]), .Z(n154) );
  AOI22M1P U170 ( .A(n56), .B(Packet_From_Link_N[30]), .C(n61), .D(
        Packet_From_Link_S[30]), .Z(n153) );
  AOI22M1P U171 ( .A(n58), .B(Packet_From_Link_W[30]), .C(n51), .D(
        Packet_From_Node_30), .Z(n152) );
  ND3M1P U172 ( .A(n154), .B(n153), .C(n152), .Z(n264) );
  AOI22M1P U173 ( .A(chosenPacket[31]), .B(n55), .C(n63), .D(
        Packet_From_Link_E[31]), .Z(n159) );
  AOI22M1P U174 ( .A(n56), .B(Packet_From_Link_N[31]), .C(n61), .D(
        Packet_From_Link_S[31]), .Z(n158) );
  AOI22M1P U175 ( .A(n58), .B(Packet_From_Link_W[31]), .C(n51), .D(
        Packet_From_Node_31), .Z(n157) );
  ND3M1P U176 ( .A(n159), .B(n158), .C(n157), .Z(n263) );
  AO21CNM1P U177 ( .A(n8), .B(n160), .C(Rst_n), .Z(n188) );
  AOI22M1P U178 ( .A(chosenPacket[23]), .B(n188), .C(N115), .D(n233), .Z(n163)
         );
  AOI22M1P U179 ( .A(n58), .B(Packet_From_Link_W[23]), .C(n56), .D(
        Packet_From_Link_N[23]), .Z(n162) );
  AOI22M1P U180 ( .A(n63), .B(Packet_From_Link_E[23]), .C(n61), .D(
        Packet_From_Link_S[23]), .Z(n161) );
  ND3M1P U181 ( .A(n163), .B(n162), .C(n161), .Z(n262) );
  N1M1P U182 ( .A(chosenPacket[24]), .Z(n238) );
  N1M1P U183 ( .A(chosenPacket[28]), .Z(n236) );
  ND2M1P U184 ( .A(Router_Address[3]), .B(n44), .Z(n212) );
  ND2M1P U185 ( .A(Router_Address[4]), .B(n236), .Z(n216) );
  OAI211M1P U186 ( .A(Router_Address[4]), .B(n236), .C(n212), .D(n216), .Z(
        n167) );
  NR2M1P U187 ( .A(Router_Address[5]), .B(n43), .Z(n215) );
  NR2M1P U188 ( .A(Router_Address[6]), .B(n42), .Z(n218) );
  NR2M1P U189 ( .A(n215), .B(n218), .Z(n222) );
  AOI22M1P U190 ( .A(Router_Address[5]), .B(n43), .C(Router_Address[6]), .D(
        n42), .Z(n214) );
  NR2M1P U191 ( .A(Router_Address[3]), .B(n44), .Z(n164) );
  NR2M1P U192 ( .A(Router_Address[0]), .B(n238), .Z(n201) );
  AOI211M1P U193 ( .A(Router_Address[1]), .B(n45), .C(n164), .D(n201), .Z(n165) );
  N1M1P U194 ( .A(chosenPacket[26]), .Z(n237) );
  ND2M1P U195 ( .A(Router_Address[2]), .B(n237), .Z(n200) );
  ND4M1P U196 ( .A(n222), .B(n214), .C(n165), .D(n200), .Z(n166) );
  AOI211M1P U197 ( .A(Router_Address[0]), .B(n238), .C(n167), .D(n166), .Z(
        n169) );
  OAI22M1P U198 ( .A(Router_Address[2]), .B(n237), .C(Router_Address[1]), .D(
        n45), .Z(n206) );
  AOI21M1P U199 ( .A(Router_Address[7]), .B(n41), .C(n206), .Z(n168) );
  OAI211M1P U200 ( .A(Router_Address[7]), .B(n41), .C(n169), .D(n168), .Z(n197) );
  NR2M1P U201 ( .A(n8), .B(n197), .Z(n307) );
  AO21CNM1P U202 ( .A(To_Node_Write), .B(n223), .C(n66), .Z(n261) );
  AOI22M1P U203 ( .A(chosenPacket[16]), .B(n188), .C(n233), .D(N108), .Z(n172)
         );
  AOI22M1P U204 ( .A(n63), .B(Packet_From_Link_E[16]), .C(n56), .D(
        Packet_From_Link_N[16]), .Z(n171) );
  AOI22M1P U205 ( .A(n58), .B(Packet_From_Link_W[16]), .C(n61), .D(
        Packet_From_Link_S[16]), .Z(n170) );
  ND3M1P U206 ( .A(n172), .B(n171), .C(n170), .Z(n260) );
  AOI22M1P U207 ( .A(chosenPacket[17]), .B(n188), .C(n233), .D(N109), .Z(n175)
         );
  AOI22M1P U208 ( .A(n58), .B(Packet_From_Link_W[17]), .C(n56), .D(
        Packet_From_Link_N[17]), .Z(n174) );
  AOI22M1P U209 ( .A(n63), .B(Packet_From_Link_E[17]), .C(n61), .D(
        Packet_From_Link_S[17]), .Z(n173) );
  ND3M1P U210 ( .A(n175), .B(n174), .C(n173), .Z(n259) );
  AOI22M1P U211 ( .A(chosenPacket[18]), .B(n188), .C(n233), .D(N110), .Z(n178)
         );
  AOI22M1P U212 ( .A(n58), .B(Packet_From_Link_W[18]), .C(n56), .D(
        Packet_From_Link_N[18]), .Z(n177) );
  AOI22M1P U213 ( .A(n63), .B(Packet_From_Link_E[18]), .C(n61), .D(
        Packet_From_Link_S[18]), .Z(n176) );
  ND3M1P U214 ( .A(n178), .B(n177), .C(n176), .Z(n258) );
  AOI22M1P U215 ( .A(chosenPacket[19]), .B(n188), .C(N111), .D(n233), .Z(n181)
         );
  AOI22M1P U216 ( .A(n58), .B(Packet_From_Link_W[19]), .C(n56), .D(
        Packet_From_Link_N[19]), .Z(n180) );
  AOI22M1P U217 ( .A(n63), .B(Packet_From_Link_E[19]), .C(n61), .D(
        Packet_From_Link_S[19]), .Z(n179) );
  ND3M1P U218 ( .A(n181), .B(n180), .C(n179), .Z(n257) );
  AOI22M1P U219 ( .A(chosenPacket[20]), .B(n188), .C(N112), .D(n233), .Z(n184)
         );
  AOI22M1P U220 ( .A(n58), .B(Packet_From_Link_W[20]), .C(n56), .D(
        Packet_From_Link_N[20]), .Z(n183) );
  AOI22M1P U221 ( .A(n63), .B(Packet_From_Link_E[20]), .C(n61), .D(
        Packet_From_Link_S[20]), .Z(n182) );
  ND3M1P U222 ( .A(n184), .B(n183), .C(n182), .Z(n256) );
  AOI22M1P U223 ( .A(chosenPacket[21]), .B(n188), .C(n233), .D(N113), .Z(n187)
         );
  AOI22M1P U224 ( .A(n50), .B(Packet_From_Link_W[21]), .C(n56), .D(
        Packet_From_Link_N[21]), .Z(n186) );
  AOI22M1P U225 ( .A(n63), .B(Packet_From_Link_E[21]), .C(n62), .D(
        Packet_From_Link_S[21]), .Z(n185) );
  ND3M1P U226 ( .A(n187), .B(n186), .C(n185), .Z(n255) );
  AOI22M1P U227 ( .A(chosenPacket[22]), .B(n188), .C(N114), .D(n233), .Z(n195)
         );
  AOI22M1P U228 ( .A(n50), .B(Packet_From_Link_W[22]), .C(n56), .D(
        Packet_From_Link_N[22]), .Z(n194) );
  AOI22M1P U229 ( .A(n63), .B(Packet_From_Link_E[22]), .C(n62), .D(
        Packet_From_Link_S[22]), .Z(n193) );
  ND3M1P U230 ( .A(n195), .B(n194), .C(n193), .Z(n254) );
  ND4M1P U231 ( .A(chosenPacket[17]), .B(chosenPacket[18]), .C(
        chosenPacket[19]), .D(N108), .Z(n199) );
  ND4M1P U232 ( .A(N115), .B(N114), .C(N112), .D(n196), .Z(n198) );
  OA21M1P U233 ( .A(n199), .B(n198), .C(n197), .Z(n205) );
  N1M1P U234 ( .A(n200), .Z(n210) );
  ND2M1P U235 ( .A(Router_Address[1]), .B(n45), .Z(n208) );
  AOI21M1P U236 ( .A(n201), .B(n208), .C(n206), .Z(n202) );
  OAI22M1P U237 ( .A(n210), .B(n202), .C(Router_Address[3]), .D(n44), .Z(n203)
         );
  ND4DNM1P U238 ( .D(TxQueue_Full_N), .A(Link_Config[3]), .B(n203), .C(n212), 
        .Z(n204) );
  NR2BNM1P U239 ( .B(n205), .A(n204), .Z(n231) );
  OA21M1P U240 ( .A(n231), .B(TxQueue_Write_N), .C(n223), .Z(n253) );
  ND2M1P U241 ( .A(n205), .B(n204), .Z(n234) );
  ND2M1P U242 ( .A(Router_Address[0]), .B(n238), .Z(n207) );
  AOI21M1P U243 ( .A(n208), .B(n207), .C(n206), .Z(n209) );
  OAI22M1P U244 ( .A(n210), .B(n209), .C(Router_Address[3]), .D(n44), .Z(n211)
         );
  AOI21M1P U245 ( .A(n212), .B(n211), .C(TxQueue_Full_S), .Z(n213) );
  ND2M1P U246 ( .A(Link_Config[2]), .B(n213), .Z(n232) );
  NR2M1P U247 ( .A(n234), .B(n232), .Z(n230) );
  OA21M1P U248 ( .A(n230), .B(TxQueue_Write_S), .C(n223), .Z(n252) );
  N1M1P U249 ( .A(Router_Address[7]), .Z(n220) );
  OAI21M1P U250 ( .A(n216), .B(n215), .C(n214), .Z(n217) );
  ND2BNM1P U251 ( .B(n218), .A(n217), .Z(n219) );
  MAJN3M1P U252 ( .A(chosenPacket[31]), .B(n220), .C(n219), .Z(n221) );
  ND3CNM1P U253 ( .C(TxQueue_Full_W), .A(Link_Config[1]), .B(n221), .Z(n303)
         );
  NR3CNM1P U254 ( .C(n232), .A(n234), .B(n8), .Z(n304) );
  N1M1P U255 ( .A(n304), .Z(n224) );
  OAI22CDNM1P U256 ( .A(n303), .B(n224), .C(n223), .D(TxQueue_Write_W), .Z(
        n251) );
  OAI22CDNM1P U257 ( .A(n302), .B(n224), .C(n223), .D(TxQueue_Write_E), .Z(
        n250) );
  N1M1P U258 ( .A(n305), .Z(n229) );
  OAI22CDNM1P U259 ( .A(n6), .B(n229), .C(n8), .D(RxQueue_Read_E), .Z(n249) );
  AOI22M1P U260 ( .A(n8), .B(RxQueue_Read_W), .C(n225), .D(n305), .Z(n226) );
  OAI22CDNM1P U261 ( .A(n227), .B(n229), .C(n8), .D(RxQueue_Read_S), .Z(n247)
         );
  OAI22CDNM1P U262 ( .A(n228), .B(n229), .C(n8), .D(RxQueue_Read_N), .Z(n246)
         );
  OAI22CDNM1P U263 ( .A(n57), .B(n229), .C(n8), .D(Node_Read), .Z(n245) );
  ND3CNM1P U264 ( .C(n234), .A(n233), .B(n232), .Z(n235) );
  NR2M1P U265 ( .A(n303), .B(n235), .Z(n38) );
  NR2M1P U266 ( .A(n302), .B(n235), .Z(n37) );
  AOI22DNM1P U267 ( .A(n65), .B(n236), .D(Packet_To_Node[28]), .C(n66), .Z(n35) );
  AOI22DNM1P U268 ( .A(n65), .B(n237), .D(Packet_To_Node[26]), .C(n66), .Z(n34) );
  AOI22DNM1P U269 ( .A(n65), .B(n238), .D(Packet_To_Node[24]), .C(n66), .Z(n33) );
  OAI22M1P U270 ( .A(n66), .B(N115), .C(Packet_To_Node[23]), .D(n65), .Z(n239)
         );
  N1M1P U271 ( .A(n239), .Z(n32) );
  AOI22DNM1P U272 ( .A(n65), .B(n240), .D(Packet_To_Node[21]), .C(n66), .Z(n30) );
  OAI22M1P U273 ( .A(n66), .B(N112), .C(Packet_To_Node[20]), .D(n65), .Z(n241)
         );
  N1M1P U274 ( .A(n241), .Z(n29) );
  AOI22DNM1P U275 ( .A(n65), .B(n242), .D(Packet_To_Node[19]), .C(n66), .Z(n28) );
  OAI22M1P U276 ( .A(n66), .B(N110), .C(Packet_To_Node[18]), .D(n65), .Z(n243)
         );
  N1M1P U277 ( .A(n243), .Z(n27) );
  AOI22DNM1P U278 ( .A(n65), .B(n244), .D(Packet_To_Node[17]), .C(n66), .Z(n26) );
  AOI22DNM1P U279 ( .A(n65), .B(chosenPacket[16]), .D(Packet_To_Node[16]), .C(
        n66), .Z(n25) );
  OAI22M1P U280 ( .A(n66), .B(chosenPacket[15]), .C(Packet_To_Node[15]), .D(
        n65), .Z(n248) );
  N1M1P U281 ( .A(n248), .Z(n24) );
  OAI22M1P U282 ( .A(n66), .B(chosenPacket[14]), .C(Packet_To_Node[14]), .D(
        n65), .Z(n287) );
  N1M1P U283 ( .A(n287), .Z(n23) );
  OAI22M1P U284 ( .A(n66), .B(chosenPacket[13]), .C(Packet_To_Node[13]), .D(
        n107), .Z(n288) );
  N1M1P U285 ( .A(n288), .Z(n22) );
  OAI22M1P U286 ( .A(n66), .B(chosenPacket[12]), .C(Packet_To_Node[12]), .D(
        n107), .Z(n289) );
  N1M1P U287 ( .A(n289), .Z(n21) );
  OAI22M1P U288 ( .A(n66), .B(chosenPacket[11]), .C(Packet_To_Node[11]), .D(
        n107), .Z(n290) );
  N1M1P U289 ( .A(n290), .Z(n20) );
  OAI22M1P U290 ( .A(n66), .B(chosenPacket[10]), .C(Packet_To_Node[10]), .D(
        n107), .Z(n291) );
  N1M1P U291 ( .A(n291), .Z(n19) );
  OAI22M1P U292 ( .A(n66), .B(chosenPacket[9]), .C(Packet_To_Node[9]), .D(n107), .Z(n292) );
  N1M1P U293 ( .A(n292), .Z(n18) );
  OAI22M1P U294 ( .A(n66), .B(chosenPacket[8]), .C(Packet_To_Node[8]), .D(n107), .Z(n293) );
  N1M1P U295 ( .A(n293), .Z(n17) );
  OAI22M1P U296 ( .A(n66), .B(chosenPacket[7]), .C(Packet_To_Node[7]), .D(n65), 
        .Z(n294) );
  N1M1P U297 ( .A(n294), .Z(n16) );
  OAI22M1P U298 ( .A(n66), .B(chosenPacket[6]), .C(Packet_To_Node[6]), .D(n65), 
        .Z(n295) );
  N1M1P U299 ( .A(n295), .Z(n15) );
  OAI22M1P U300 ( .A(n66), .B(chosenPacket[5]), .C(Packet_To_Node[5]), .D(n65), 
        .Z(n296) );
  N1M1P U301 ( .A(n296), .Z(n14) );
  OAI22M1P U302 ( .A(n66), .B(chosenPacket[4]), .C(Packet_To_Node[4]), .D(n65), 
        .Z(n297) );
  N1M1P U303 ( .A(n297), .Z(n13) );
  OAI22M1P U304 ( .A(n66), .B(chosenPacket[3]), .C(Packet_To_Node[3]), .D(n65), 
        .Z(n298) );
  N1M1P U305 ( .A(n298), .Z(n12) );
  OAI22M1P U306 ( .A(n66), .B(chosenPacket[2]), .C(Packet_To_Node[2]), .D(n65), 
        .Z(n299) );
  N1M1P U307 ( .A(n299), .Z(n11) );
  OAI22M1P U308 ( .A(n66), .B(chosenPacket[1]), .C(Packet_To_Node[1]), .D(n65), 
        .Z(n300) );
  N1M1P U309 ( .A(n300), .Z(n10) );
  OAI22M1P U310 ( .A(n66), .B(chosenPacket[0]), .C(Packet_To_Node[0]), .D(n65), 
        .Z(n301) );
  N1M1P U311 ( .A(n301), .Z(n9) );
  AND3M1P U312 ( .A(n304), .B(n303), .C(n302), .Z(n306) );
  AOI211M1P U313 ( .A(To_Node_Full), .B(n307), .C(n306), .D(n305), .Z(n7) );
  N1M1P U314 ( .A(n5), .Z(Packet_To_Node[31]) );
  N1M1P U315 ( .A(n4), .Z(Packet_To_Node[30]) );
  N1M1P U316 ( .A(n3), .Z(Packet_To_Node[29]) );
  N1M1P U317 ( .A(n2), .Z(Packet_To_Node[27]) );
  N1M1P U318 ( .A(n1), .Z(Packet_To_Node[25]) );
endmodule


module Packet_Queue_1 ( Clk_r, Rst_n, Packet_In, Read_Ack, Write_Ack, 
        Packet_Out, Empty, Full );
  input [31:0] Packet_In;
  output [31:0] Packet_Out;
  input Clk_r, Rst_n, Read_Ack, Write_Ack;
  output Empty, Full;
  wire   \Queue[4][31] , \Queue[4][30] , \Queue[4][29] , \Queue[4][28] ,
         \Queue[4][27] , \Queue[4][26] , \Queue[4][25] , \Queue[4][24] ,
         \Queue[4][23] , \Queue[4][22] , \Queue[4][21] , \Queue[4][20] ,
         \Queue[4][19] , \Queue[4][18] , \Queue[4][17] , \Queue[4][16] ,
         \Queue[4][15] , \Queue[4][14] , \Queue[4][13] , \Queue[4][12] ,
         \Queue[4][11] , \Queue[4][10] , \Queue[4][9] , \Queue[4][8] ,
         \Queue[4][7] , \Queue[4][6] , \Queue[4][5] , \Queue[4][4] ,
         \Queue[4][3] , \Queue[4][2] , \Queue[4][1] , \Queue[4][0] ,
         \Queue[3][31] , \Queue[3][30] , \Queue[3][29] , \Queue[3][28] ,
         \Queue[3][27] , \Queue[3][26] , \Queue[3][25] , \Queue[3][24] ,
         \Queue[3][23] , \Queue[3][22] , \Queue[3][21] , \Queue[3][20] ,
         \Queue[3][19] , \Queue[3][18] , \Queue[3][17] , \Queue[3][16] ,
         \Queue[3][15] , \Queue[3][14] , \Queue[3][13] , \Queue[3][12] ,
         \Queue[3][11] , \Queue[3][10] , \Queue[3][9] , \Queue[3][8] ,
         \Queue[3][7] , \Queue[3][6] , \Queue[3][5] , \Queue[3][4] ,
         \Queue[3][3] , \Queue[3][2] , \Queue[3][1] , \Queue[3][0] ,
         \Queue[2][31] , \Queue[2][30] , \Queue[2][29] , \Queue[2][28] ,
         \Queue[2][27] , \Queue[2][26] , \Queue[2][25] , \Queue[2][24] ,
         \Queue[2][23] , \Queue[2][22] , \Queue[2][21] , \Queue[2][20] ,
         \Queue[2][19] , \Queue[2][18] , \Queue[2][17] , \Queue[2][16] ,
         \Queue[2][15] , \Queue[2][14] , \Queue[2][13] , \Queue[2][12] ,
         \Queue[2][11] , \Queue[2][10] , \Queue[2][9] , \Queue[2][8] ,
         \Queue[2][7] , \Queue[2][6] , \Queue[2][5] , \Queue[2][4] ,
         \Queue[2][3] , \Queue[2][2] , \Queue[2][1] , \Queue[2][0] ,
         \Queue[1][31] , \Queue[1][30] , \Queue[1][29] , \Queue[1][28] ,
         \Queue[1][27] , \Queue[1][26] , \Queue[1][25] , \Queue[1][24] ,
         \Queue[1][23] , \Queue[1][22] , \Queue[1][21] , \Queue[1][20] ,
         \Queue[1][19] , \Queue[1][18] , \Queue[1][17] , \Queue[1][16] ,
         \Queue[1][15] , \Queue[1][14] , \Queue[1][13] , \Queue[1][12] ,
         \Queue[1][11] , \Queue[1][10] , \Queue[1][9] , \Queue[1][8] ,
         \Queue[1][7] , \Queue[1][6] , \Queue[1][5] , \Queue[1][4] ,
         \Queue[1][3] , \Queue[1][2] , \Queue[1][1] , \Queue[1][0] , n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549;
  wire   [2:0] Count;

  FDN2QM1P \Count_reg[0]  ( .D(n384), .CPN(Clk_r), .CD(n19), .Q(Count[0]) );
  FDN2QM1P \Count_reg[1]  ( .D(n385), .CPN(Clk_r), .CD(n19), .Q(Count[1]) );
  FDN2QM1P \Count_reg[2]  ( .D(n386), .CPN(Clk_r), .CD(n19), .Q(Count[2]) );
  FDN1QM1P \Queue_reg[4][30]  ( .D(n418), .CPN(Clk_r), .Q(\Queue[4][30] ) );
  FDN1QM1P \Queue_reg[3][30]  ( .D(n546), .CPN(Clk_r), .Q(\Queue[3][30] ) );
  FDN1QM1P \Queue_reg[2][30]  ( .D(n514), .CPN(Clk_r), .Q(\Queue[2][30] ) );
  FDN1QM1P \Queue_reg[4][29]  ( .D(n417), .CPN(Clk_r), .Q(\Queue[4][29] ) );
  FDN1QM1P \Queue_reg[3][29]  ( .D(n545), .CPN(Clk_r), .Q(\Queue[3][29] ) );
  FDN1QM1P \Queue_reg[2][29]  ( .D(n513), .CPN(Clk_r), .Q(\Queue[2][29] ) );
  FDN1QM1P \Queue_reg[4][28]  ( .D(n416), .CPN(Clk_r), .Q(\Queue[4][28] ) );
  FDN1QM1P \Queue_reg[3][28]  ( .D(n544), .CPN(Clk_r), .Q(\Queue[3][28] ) );
  FDN1QM1P \Queue_reg[2][28]  ( .D(n512), .CPN(Clk_r), .Q(\Queue[2][28] ) );
  FDN1QM1P \Queue_reg[4][27]  ( .D(n415), .CPN(Clk_r), .Q(\Queue[4][27] ) );
  FDN1QM1P \Queue_reg[3][27]  ( .D(n543), .CPN(Clk_r), .Q(\Queue[3][27] ) );
  FDN1QM1P \Queue_reg[2][27]  ( .D(n511), .CPN(Clk_r), .Q(\Queue[2][27] ) );
  FDN1QM1P \Queue_reg[4][26]  ( .D(n414), .CPN(Clk_r), .Q(\Queue[4][26] ) );
  FDN1QM1P \Queue_reg[3][26]  ( .D(n542), .CPN(Clk_r), .Q(\Queue[3][26] ) );
  FDN1QM1P \Queue_reg[2][26]  ( .D(n510), .CPN(Clk_r), .Q(\Queue[2][26] ) );
  FDN1QM1P \Queue_reg[4][25]  ( .D(n413), .CPN(Clk_r), .Q(\Queue[4][25] ) );
  FDN1QM1P \Queue_reg[3][25]  ( .D(n541), .CPN(Clk_r), .Q(\Queue[3][25] ) );
  FDN1QM1P \Queue_reg[2][25]  ( .D(n509), .CPN(Clk_r), .Q(\Queue[2][25] ) );
  FDN1QM1P \Queue_reg[4][24]  ( .D(n412), .CPN(Clk_r), .Q(\Queue[4][24] ) );
  FDN1QM1P \Queue_reg[3][24]  ( .D(n540), .CPN(Clk_r), .Q(\Queue[3][24] ) );
  FDN1QM1P \Queue_reg[2][24]  ( .D(n508), .CPN(Clk_r), .Q(\Queue[2][24] ) );
  FDN1QM1P \Queue_reg[4][23]  ( .D(n411), .CPN(Clk_r), .Q(\Queue[4][23] ) );
  FDN1QM1P \Queue_reg[3][23]  ( .D(n539), .CPN(Clk_r), .Q(\Queue[3][23] ) );
  FDN1QM1P \Queue_reg[2][23]  ( .D(n507), .CPN(Clk_r), .Q(\Queue[2][23] ) );
  FDN1QM1P \Queue_reg[4][22]  ( .D(n410), .CPN(Clk_r), .Q(\Queue[4][22] ) );
  FDN1QM1P \Queue_reg[3][22]  ( .D(n538), .CPN(Clk_r), .Q(\Queue[3][22] ) );
  FDN1QM1P \Queue_reg[2][22]  ( .D(n506), .CPN(Clk_r), .Q(\Queue[2][22] ) );
  FDN1QM1P \Queue_reg[4][21]  ( .D(n409), .CPN(Clk_r), .Q(\Queue[4][21] ) );
  FDN1QM1P \Queue_reg[3][21]  ( .D(n537), .CPN(Clk_r), .Q(\Queue[3][21] ) );
  FDN1QM1P \Queue_reg[2][21]  ( .D(n505), .CPN(Clk_r), .Q(\Queue[2][21] ) );
  FDN1QM1P \Queue_reg[4][20]  ( .D(n408), .CPN(Clk_r), .Q(\Queue[4][20] ) );
  FDN1QM1P \Queue_reg[3][20]  ( .D(n536), .CPN(Clk_r), .Q(\Queue[3][20] ) );
  FDN1QM1P \Queue_reg[2][20]  ( .D(n504), .CPN(Clk_r), .Q(\Queue[2][20] ) );
  FDN1QM1P \Queue_reg[4][19]  ( .D(n407), .CPN(Clk_r), .Q(\Queue[4][19] ) );
  FDN1QM1P \Queue_reg[3][19]  ( .D(n535), .CPN(Clk_r), .Q(\Queue[3][19] ) );
  FDN1QM1P \Queue_reg[2][19]  ( .D(n503), .CPN(Clk_r), .Q(\Queue[2][19] ) );
  FDN1QM1P \Queue_reg[4][18]  ( .D(n406), .CPN(Clk_r), .Q(\Queue[4][18] ) );
  FDN1QM1P \Queue_reg[3][18]  ( .D(n534), .CPN(Clk_r), .Q(\Queue[3][18] ) );
  FDN1QM1P \Queue_reg[2][18]  ( .D(n502), .CPN(Clk_r), .Q(\Queue[2][18] ) );
  FDN1QM1P \Queue_reg[4][17]  ( .D(n405), .CPN(Clk_r), .Q(\Queue[4][17] ) );
  FDN1QM1P \Queue_reg[3][17]  ( .D(n533), .CPN(Clk_r), .Q(\Queue[3][17] ) );
  FDN1QM1P \Queue_reg[2][17]  ( .D(n501), .CPN(Clk_r), .Q(\Queue[2][17] ) );
  FDN1QM1P \Queue_reg[4][16]  ( .D(n404), .CPN(Clk_r), .Q(\Queue[4][16] ) );
  FDN1QM1P \Queue_reg[3][16]  ( .D(n532), .CPN(Clk_r), .Q(\Queue[3][16] ) );
  FDN1QM1P \Queue_reg[2][16]  ( .D(n500), .CPN(Clk_r), .Q(\Queue[2][16] ) );
  FDN1QM1P \Queue_reg[4][15]  ( .D(n403), .CPN(Clk_r), .Q(\Queue[4][15] ) );
  FDN1QM1P \Queue_reg[3][15]  ( .D(n531), .CPN(Clk_r), .Q(\Queue[3][15] ) );
  FDN1QM1P \Queue_reg[2][15]  ( .D(n499), .CPN(Clk_r), .Q(\Queue[2][15] ) );
  FDN1QM1P \Queue_reg[4][14]  ( .D(n402), .CPN(Clk_r), .Q(\Queue[4][14] ) );
  FDN1QM1P \Queue_reg[3][14]  ( .D(n530), .CPN(Clk_r), .Q(\Queue[3][14] ) );
  FDN1QM1P \Queue_reg[2][14]  ( .D(n498), .CPN(Clk_r), .Q(\Queue[2][14] ) );
  FDN1QM1P \Queue_reg[4][13]  ( .D(n401), .CPN(Clk_r), .Q(\Queue[4][13] ) );
  FDN1QM1P \Queue_reg[3][13]  ( .D(n529), .CPN(Clk_r), .Q(\Queue[3][13] ) );
  FDN1QM1P \Queue_reg[2][13]  ( .D(n497), .CPN(Clk_r), .Q(\Queue[2][13] ) );
  FDN1QM1P \Queue_reg[4][12]  ( .D(n400), .CPN(Clk_r), .Q(\Queue[4][12] ) );
  FDN1QM1P \Queue_reg[3][12]  ( .D(n528), .CPN(Clk_r), .Q(\Queue[3][12] ) );
  FDN1QM1P \Queue_reg[2][12]  ( .D(n496), .CPN(Clk_r), .Q(\Queue[2][12] ) );
  FDN1QM1P \Queue_reg[4][11]  ( .D(n399), .CPN(Clk_r), .Q(\Queue[4][11] ) );
  FDN1QM1P \Queue_reg[3][11]  ( .D(n527), .CPN(Clk_r), .Q(\Queue[3][11] ) );
  FDN1QM1P \Queue_reg[2][11]  ( .D(n495), .CPN(Clk_r), .Q(\Queue[2][11] ) );
  FDN1QM1P \Queue_reg[4][10]  ( .D(n398), .CPN(Clk_r), .Q(\Queue[4][10] ) );
  FDN1QM1P \Queue_reg[3][10]  ( .D(n526), .CPN(Clk_r), .Q(\Queue[3][10] ) );
  FDN1QM1P \Queue_reg[2][10]  ( .D(n494), .CPN(Clk_r), .Q(\Queue[2][10] ) );
  FDN1QM1P \Queue_reg[4][9]  ( .D(n397), .CPN(Clk_r), .Q(\Queue[4][9] ) );
  FDN1QM1P \Queue_reg[3][9]  ( .D(n525), .CPN(Clk_r), .Q(\Queue[3][9] ) );
  FDN1QM1P \Queue_reg[2][9]  ( .D(n493), .CPN(Clk_r), .Q(\Queue[2][9] ) );
  FDN1QM1P \Queue_reg[4][8]  ( .D(n396), .CPN(Clk_r), .Q(\Queue[4][8] ) );
  FDN1QM1P \Queue_reg[3][8]  ( .D(n524), .CPN(Clk_r), .Q(\Queue[3][8] ) );
  FDN1QM1P \Queue_reg[2][8]  ( .D(n492), .CPN(Clk_r), .Q(\Queue[2][8] ) );
  FDN1QM1P \Queue_reg[4][7]  ( .D(n395), .CPN(Clk_r), .Q(\Queue[4][7] ) );
  FDN1QM1P \Queue_reg[3][7]  ( .D(n523), .CPN(Clk_r), .Q(\Queue[3][7] ) );
  FDN1QM1P \Queue_reg[2][7]  ( .D(n491), .CPN(Clk_r), .Q(\Queue[2][7] ) );
  FDN1QM1P \Queue_reg[4][6]  ( .D(n394), .CPN(Clk_r), .Q(\Queue[4][6] ) );
  FDN1QM1P \Queue_reg[3][6]  ( .D(n522), .CPN(Clk_r), .Q(\Queue[3][6] ) );
  FDN1QM1P \Queue_reg[2][6]  ( .D(n490), .CPN(Clk_r), .Q(\Queue[2][6] ) );
  FDN1QM1P \Queue_reg[4][5]  ( .D(n393), .CPN(Clk_r), .Q(\Queue[4][5] ) );
  FDN1QM1P \Queue_reg[3][5]  ( .D(n521), .CPN(Clk_r), .Q(\Queue[3][5] ) );
  FDN1QM1P \Queue_reg[2][5]  ( .D(n489), .CPN(Clk_r), .Q(\Queue[2][5] ) );
  FDN1QM1P \Queue_reg[4][4]  ( .D(n392), .CPN(Clk_r), .Q(\Queue[4][4] ) );
  FDN1QM1P \Queue_reg[3][4]  ( .D(n520), .CPN(Clk_r), .Q(\Queue[3][4] ) );
  FDN1QM1P \Queue_reg[2][4]  ( .D(n488), .CPN(Clk_r), .Q(\Queue[2][4] ) );
  FDN1QM1P \Queue_reg[4][3]  ( .D(n391), .CPN(Clk_r), .Q(\Queue[4][3] ) );
  FDN1QM1P \Queue_reg[3][3]  ( .D(n519), .CPN(Clk_r), .Q(\Queue[3][3] ) );
  FDN1QM1P \Queue_reg[2][3]  ( .D(n487), .CPN(Clk_r), .Q(\Queue[2][3] ) );
  FDN1QM1P \Queue_reg[4][2]  ( .D(n390), .CPN(Clk_r), .Q(\Queue[4][2] ) );
  FDN1QM1P \Queue_reg[3][2]  ( .D(n518), .CPN(Clk_r), .Q(\Queue[3][2] ) );
  FDN1QM1P \Queue_reg[2][2]  ( .D(n486), .CPN(Clk_r), .Q(\Queue[2][2] ) );
  FDN1QM1P \Queue_reg[4][1]  ( .D(n389), .CPN(Clk_r), .Q(\Queue[4][1] ) );
  FDN1QM1P \Queue_reg[3][1]  ( .D(n517), .CPN(Clk_r), .Q(\Queue[3][1] ) );
  FDN1QM1P \Queue_reg[2][1]  ( .D(n485), .CPN(Clk_r), .Q(\Queue[2][1] ) );
  FDN1QM1P \Queue_reg[4][0]  ( .D(n388), .CPN(Clk_r), .Q(\Queue[4][0] ) );
  FDN1QM1P \Queue_reg[3][0]  ( .D(n516), .CPN(Clk_r), .Q(\Queue[3][0] ) );
  FDN1QM1P \Queue_reg[2][0]  ( .D(n484), .CPN(Clk_r), .Q(\Queue[2][0] ) );
  FDN1QM1P \Queue_reg[4][31]  ( .D(n387), .CPN(Clk_r), .Q(\Queue[4][31] ) );
  FDN1QM1P \Queue_reg[3][31]  ( .D(n547), .CPN(Clk_r), .Q(\Queue[3][31] ) );
  FDN1QM1P \Queue_reg[2][31]  ( .D(n515), .CPN(Clk_r), .Q(\Queue[2][31] ) );
  FDN2QM1P Full_reg ( .D(n419), .CPN(Clk_r), .CD(n19), .Q(Full) );
  FDN1QM1P \Queue_reg[1][31]  ( .D(n451), .CPN(Clk_r), .Q(\Queue[1][31] ) );
  FDN1QM1P \Queue_reg[0][31]  ( .D(n483), .CPN(Clk_r), .Q(Packet_Out[31]) );
  FDN1QM1P \Queue_reg[1][30]  ( .D(n450), .CPN(Clk_r), .Q(\Queue[1][30] ) );
  FDN1QM1P \Queue_reg[0][30]  ( .D(n482), .CPN(Clk_r), .Q(Packet_Out[30]) );
  FDN1QM1P \Queue_reg[1][29]  ( .D(n449), .CPN(Clk_r), .Q(\Queue[1][29] ) );
  FDN1QM1P \Queue_reg[0][29]  ( .D(n481), .CPN(Clk_r), .Q(Packet_Out[29]) );
  FDN1QM1P \Queue_reg[1][28]  ( .D(n448), .CPN(Clk_r), .Q(\Queue[1][28] ) );
  FDN1QM1P \Queue_reg[0][28]  ( .D(n480), .CPN(Clk_r), .Q(Packet_Out[28]) );
  FDN1QM1P \Queue_reg[1][27]  ( .D(n447), .CPN(Clk_r), .Q(\Queue[1][27] ) );
  FDN1QM1P \Queue_reg[0][27]  ( .D(n479), .CPN(Clk_r), .Q(Packet_Out[27]) );
  FDN1QM1P \Queue_reg[1][26]  ( .D(n446), .CPN(Clk_r), .Q(\Queue[1][26] ) );
  FDN1QM1P \Queue_reg[0][26]  ( .D(n478), .CPN(Clk_r), .Q(Packet_Out[26]) );
  FDN1QM1P \Queue_reg[1][25]  ( .D(n445), .CPN(Clk_r), .Q(\Queue[1][25] ) );
  FDN1QM1P \Queue_reg[0][25]  ( .D(n477), .CPN(Clk_r), .Q(Packet_Out[25]) );
  FDN1QM1P \Queue_reg[1][24]  ( .D(n444), .CPN(Clk_r), .Q(\Queue[1][24] ) );
  FDN1QM1P \Queue_reg[0][24]  ( .D(n476), .CPN(Clk_r), .Q(Packet_Out[24]) );
  FDN1QM1P \Queue_reg[1][23]  ( .D(n443), .CPN(Clk_r), .Q(\Queue[1][23] ) );
  FDN1QM1P \Queue_reg[0][23]  ( .D(n475), .CPN(Clk_r), .Q(Packet_Out[23]) );
  FDN1QM1P \Queue_reg[1][22]  ( .D(n442), .CPN(Clk_r), .Q(\Queue[1][22] ) );
  FDN1QM1P \Queue_reg[0][22]  ( .D(n474), .CPN(Clk_r), .Q(Packet_Out[22]) );
  FDN1QM1P \Queue_reg[1][21]  ( .D(n441), .CPN(Clk_r), .Q(\Queue[1][21] ) );
  FDN1QM1P \Queue_reg[0][21]  ( .D(n473), .CPN(Clk_r), .Q(Packet_Out[21]) );
  FDN1QM1P \Queue_reg[1][20]  ( .D(n440), .CPN(Clk_r), .Q(\Queue[1][20] ) );
  FDN1QM1P \Queue_reg[0][20]  ( .D(n472), .CPN(Clk_r), .Q(Packet_Out[20]) );
  FDN1QM1P \Queue_reg[1][19]  ( .D(n439), .CPN(Clk_r), .Q(\Queue[1][19] ) );
  FDN1QM1P \Queue_reg[0][19]  ( .D(n471), .CPN(Clk_r), .Q(Packet_Out[19]) );
  FDN1QM1P \Queue_reg[1][18]  ( .D(n438), .CPN(Clk_r), .Q(\Queue[1][18] ) );
  FDN1QM1P \Queue_reg[0][18]  ( .D(n470), .CPN(Clk_r), .Q(Packet_Out[18]) );
  FDN1QM1P \Queue_reg[1][17]  ( .D(n437), .CPN(Clk_r), .Q(\Queue[1][17] ) );
  FDN1QM1P \Queue_reg[0][17]  ( .D(n469), .CPN(Clk_r), .Q(Packet_Out[17]) );
  FDN1QM1P \Queue_reg[1][16]  ( .D(n436), .CPN(Clk_r), .Q(\Queue[1][16] ) );
  FDN1QM1P \Queue_reg[0][16]  ( .D(n468), .CPN(Clk_r), .Q(Packet_Out[16]) );
  FDN1QM1P \Queue_reg[1][15]  ( .D(n435), .CPN(Clk_r), .Q(\Queue[1][15] ) );
  FDN1QM1P \Queue_reg[0][15]  ( .D(n467), .CPN(Clk_r), .Q(Packet_Out[15]) );
  FDN1QM1P \Queue_reg[1][14]  ( .D(n434), .CPN(Clk_r), .Q(\Queue[1][14] ) );
  FDN1QM1P \Queue_reg[0][14]  ( .D(n466), .CPN(Clk_r), .Q(Packet_Out[14]) );
  FDN1QM1P \Queue_reg[1][13]  ( .D(n433), .CPN(Clk_r), .Q(\Queue[1][13] ) );
  FDN1QM1P \Queue_reg[0][13]  ( .D(n465), .CPN(Clk_r), .Q(Packet_Out[13]) );
  FDN1QM1P \Queue_reg[1][12]  ( .D(n432), .CPN(Clk_r), .Q(\Queue[1][12] ) );
  FDN1QM1P \Queue_reg[0][12]  ( .D(n464), .CPN(Clk_r), .Q(Packet_Out[12]) );
  FDN1QM1P \Queue_reg[1][11]  ( .D(n431), .CPN(Clk_r), .Q(\Queue[1][11] ) );
  FDN1QM1P \Queue_reg[0][11]  ( .D(n463), .CPN(Clk_r), .Q(Packet_Out[11]) );
  FDN1QM1P \Queue_reg[1][10]  ( .D(n430), .CPN(Clk_r), .Q(\Queue[1][10] ) );
  FDN1QM1P \Queue_reg[0][10]  ( .D(n462), .CPN(Clk_r), .Q(Packet_Out[10]) );
  FDN1QM1P \Queue_reg[1][9]  ( .D(n429), .CPN(Clk_r), .Q(\Queue[1][9] ) );
  FDN1QM1P \Queue_reg[0][9]  ( .D(n461), .CPN(Clk_r), .Q(Packet_Out[9]) );
  FDN1QM1P \Queue_reg[1][8]  ( .D(n428), .CPN(Clk_r), .Q(\Queue[1][8] ) );
  FDN1QM1P \Queue_reg[0][8]  ( .D(n460), .CPN(Clk_r), .Q(Packet_Out[8]) );
  FDN1QM1P \Queue_reg[1][7]  ( .D(n427), .CPN(Clk_r), .Q(\Queue[1][7] ) );
  FDN1QM1P \Queue_reg[0][7]  ( .D(n459), .CPN(Clk_r), .Q(Packet_Out[7]) );
  FDN1QM1P \Queue_reg[1][6]  ( .D(n426), .CPN(Clk_r), .Q(\Queue[1][6] ) );
  FDN1QM1P \Queue_reg[0][6]  ( .D(n458), .CPN(Clk_r), .Q(Packet_Out[6]) );
  FDN1QM1P \Queue_reg[1][5]  ( .D(n425), .CPN(Clk_r), .Q(\Queue[1][5] ) );
  FDN1QM1P \Queue_reg[0][5]  ( .D(n457), .CPN(Clk_r), .Q(Packet_Out[5]) );
  FDN1QM1P \Queue_reg[1][4]  ( .D(n424), .CPN(Clk_r), .Q(\Queue[1][4] ) );
  FDN1QM1P \Queue_reg[0][4]  ( .D(n456), .CPN(Clk_r), .Q(Packet_Out[4]) );
  FDN1QM1P \Queue_reg[1][3]  ( .D(n423), .CPN(Clk_r), .Q(\Queue[1][3] ) );
  FDN1QM1P \Queue_reg[0][3]  ( .D(n455), .CPN(Clk_r), .Q(Packet_Out[3]) );
  FDN1QM1P \Queue_reg[1][2]  ( .D(n422), .CPN(Clk_r), .Q(\Queue[1][2] ) );
  FDN1QM1P \Queue_reg[0][2]  ( .D(n454), .CPN(Clk_r), .Q(Packet_Out[2]) );
  FDN1QM1P \Queue_reg[1][1]  ( .D(n421), .CPN(Clk_r), .Q(\Queue[1][1] ) );
  FDN1QM1P \Queue_reg[0][1]  ( .D(n453), .CPN(Clk_r), .Q(Packet_Out[1]) );
  FDN1QM1P \Queue_reg[1][0]  ( .D(n420), .CPN(Clk_r), .Q(\Queue[1][0] ) );
  FDN1QM1P \Queue_reg[0][0]  ( .D(n452), .CPN(Clk_r), .Q(Packet_Out[0]) );
  FDN2QM1P Empty_reg ( .D(n549), .CPN(Clk_r), .CD(n19), .Q(n548) );
  BUFM2P U3 ( .A(n102), .Z(n5) );
  BUFM1P U4 ( .A(n101), .Z(n11) );
  BUFM2P U5 ( .A(n104), .Z(n13) );
  BUFM1P U6 ( .A(n101), .Z(n12) );
  BUFM2P U7 ( .A(n104), .Z(n14) );
  BUFM2P U8 ( .A(n139), .Z(n4) );
  BUFM2P U9 ( .A(n376), .Z(n3) );
  N1M1P U10 ( .A(Read_Ack), .Z(n144) );
  OAI211M1P U11 ( .A(n149), .B(n144), .C(n6), .D(n143), .Z(n379) );
  OAI211M1P U12 ( .A(n147), .B(n144), .C(n6), .D(n105), .Z(n142) );
  AOI21M1P U13 ( .A(n6), .B(n107), .C(n148), .Z(n64) );
  ND2M1P U14 ( .A(Read_Ack), .B(n19), .Z(n148) );
  NR2I1M8P U15 ( .A(n68), .B(n28), .Z(n27) );
  OAI211M4P U16 ( .A(n107), .B(n144), .C(n6), .D(n31), .Z(n66) );
  OAI211M4P U17 ( .A(n107), .B(n146), .C(n19), .D(n145), .Z(n140) );
  OAI21M2P U18 ( .A(n6), .B(Read_Ack), .C(n31), .Z(n63) );
  NR3M1P U19 ( .A(Count[2]), .B(n30), .C(n29), .Z(n147) );
  BUFM2P U20 ( .A(n142), .Z(n16) );
  BUFM2P U21 ( .A(n379), .Z(n18) );
  BUFM2P U22 ( .A(n142), .Z(n15) );
  BUFM2P U23 ( .A(n379), .Z(n17) );
  ND2M1P U24 ( .A(n25), .B(n19), .Z(n68) );
  N1M1P U25 ( .A(n149), .Z(n28) );
  NR2M2P U26 ( .A(Read_Ack), .B(n106), .Z(n25) );
  NR3M1P U27 ( .A(Count[0]), .B(Count[2]), .C(n29), .Z(n107) );
  NR3M1P U28 ( .A(Count[0]), .B(Count[1]), .C(n26), .Z(n149) );
  N1M3P U29 ( .A(n6), .Z(n106) );
  NR3M1P U30 ( .A(n30), .B(Count[2]), .C(Count[1]), .Z(n383) );
  N1M1P U31 ( .A(Count[0]), .Z(n30) );
  BUFM8P U32 ( .A(Write_Ack), .Z(n6) );
  N1M1P U33 ( .A(Count[1]), .Z(n29) );
  N1M1P U34 ( .A(Count[2]), .Z(n26) );
  BUFM2P U35 ( .A(Rst_n), .Z(n19) );
  OAI211M6P U36 ( .A(n383), .B(n144), .C(n6), .D(n69), .Z(n104) );
  OAI211M4P U37 ( .A(n147), .B(n146), .C(n19), .D(n145), .Z(n377) );
  N1M1P U38 ( .A(Packet_In[27]), .Z(n205) );
  N1M1P U39 ( .A(Packet_In[29]), .Z(n373) );
  N1M1P U40 ( .A(Packet_In[31]), .Z(n380) );
  N1M1P U41 ( .A(Packet_In[30]), .Z(n375) );
  N1M1P U42 ( .A(Packet_In[0]), .Z(n151) );
  N1M1P U43 ( .A(Packet_In[3]), .Z(n157) );
  N1M1P U44 ( .A(Packet_In[22]), .Z(n195) );
  N1M1P U45 ( .A(Packet_In[2]), .Z(n155) );
  N1M1P U46 ( .A(Packet_In[6]), .Z(n163) );
  N1M1P U47 ( .A(Packet_In[4]), .Z(n159) );
  N1M1P U48 ( .A(Packet_In[7]), .Z(n165) );
  N1M1P U49 ( .A(Packet_In[5]), .Z(n161) );
  N1M1P U50 ( .A(Packet_In[9]), .Z(n169) );
  N1M1P U51 ( .A(Packet_In[11]), .Z(n173) );
  N1M1P U52 ( .A(Packet_In[10]), .Z(n171) );
  N1M1P U53 ( .A(Packet_In[8]), .Z(n167) );
  N1M1P U54 ( .A(Packet_In[15]), .Z(n181) );
  N1M1P U55 ( .A(Packet_In[25]), .Z(n201) );
  N1M1P U56 ( .A(Packet_In[1]), .Z(n153) );
  N1M1P U57 ( .A(Packet_In[14]), .Z(n179) );
  N1M1P U58 ( .A(Packet_In[20]), .Z(n191) );
  N1M1P U59 ( .A(Packet_In[18]), .Z(n187) );
  N1M1P U60 ( .A(Packet_In[13]), .Z(n177) );
  N1M1P U61 ( .A(Packet_In[12]), .Z(n175) );
  N1M1P U62 ( .A(Packet_In[23]), .Z(n197) );
  N1M2P U63 ( .A(n69), .Z(n101) );
  BUFM2P U64 ( .A(n64), .Z(n10) );
  BUFM2P U65 ( .A(n63), .Z(n7) );
  BUFM2P U66 ( .A(n63), .Z(n8) );
  BUFM2P U67 ( .A(n64), .Z(n9) );
  N1M2P U68 ( .A(n25), .Z(n146) );
  NR2M1P U69 ( .A(n144), .B(n6), .Z(n382) );
  NR2M1P U70 ( .A(n25), .B(n382), .Z(n381) );
  AOI22CDNM1P U71 ( .A(n381), .B(n30), .C(n381), .D(n30), .Z(n384) );
  N1M1P U72 ( .A(n382), .Z(n24) );
  AOI22M1P U73 ( .A(Count[0]), .B(n146), .C(n24), .D(n30), .Z(n21) );
  AOI22CDNM1P U74 ( .A(Count[1]), .B(n21), .C(n21), .D(Count[1]), .Z(n385) );
  ND3M1P U75 ( .A(n30), .B(n26), .C(n29), .Z(n67) );
  ND2M1P U76 ( .A(Count[1]), .B(Read_Ack), .Z(n20) );
  OAI211M1P U77 ( .A(Count[1]), .B(n146), .C(n21), .D(n20), .Z(n22) );
  AOI22M1P U78 ( .A(n25), .B(n147), .C(Count[2]), .D(n22), .Z(n23) );
  OAI21M1P U79 ( .A(n67), .B(n24), .C(n23), .Z(n386) );
  AOI22CDNM1P U80 ( .A(n27), .B(n380), .C(\Queue[4][31] ), .D(n27), .Z(n387)
         );
  AOI22CDNM1P U81 ( .A(n27), .B(n151), .C(\Queue[4][0] ), .D(n27), .Z(n388) );
  AOI22CDNM1P U82 ( .A(n27), .B(n153), .C(\Queue[4][1] ), .D(n27), .Z(n389) );
  AOI22CDNM1P U83 ( .A(n27), .B(n155), .C(\Queue[4][2] ), .D(n27), .Z(n390) );
  AOI22CDNM1P U84 ( .A(n27), .B(n157), .C(\Queue[4][3] ), .D(n27), .Z(n391) );
  AOI22CDNM1P U85 ( .A(n27), .B(n159), .C(\Queue[4][4] ), .D(n27), .Z(n392) );
  AOI22CDNM1P U86 ( .A(n27), .B(n161), .C(\Queue[4][5] ), .D(n27), .Z(n393) );
  AOI22CDNM1P U87 ( .A(n27), .B(n163), .C(\Queue[4][6] ), .D(n27), .Z(n394) );
  AOI22CDNM1P U88 ( .A(n27), .B(n165), .C(\Queue[4][7] ), .D(n27), .Z(n395) );
  AOI22CDNM1P U89 ( .A(n27), .B(n167), .C(\Queue[4][8] ), .D(n27), .Z(n396) );
  AOI22CDNM1P U90 ( .A(n27), .B(n169), .C(\Queue[4][9] ), .D(n27), .Z(n397) );
  AOI22CDNM1P U91 ( .A(n27), .B(n171), .C(\Queue[4][10] ), .D(n27), .Z(n398)
         );
  AOI22CDNM1P U92 ( .A(n27), .B(n173), .C(\Queue[4][11] ), .D(n27), .Z(n399)
         );
  AOI22CDNM1P U93 ( .A(n27), .B(n175), .C(\Queue[4][12] ), .D(n27), .Z(n400)
         );
  AOI22CDNM1P U94 ( .A(n27), .B(n177), .C(\Queue[4][13] ), .D(n27), .Z(n401)
         );
  AOI22CDNM1P U95 ( .A(n27), .B(n179), .C(\Queue[4][14] ), .D(n27), .Z(n402)
         );
  AOI22CDNM1P U96 ( .A(n27), .B(n181), .C(\Queue[4][15] ), .D(n27), .Z(n403)
         );
  N1M1P U97 ( .A(Packet_In[16]), .Z(n183) );
  AOI22CDNM1P U98 ( .A(n27), .B(n183), .C(\Queue[4][16] ), .D(n27), .Z(n404)
         );
  N1M1P U99 ( .A(Packet_In[17]), .Z(n185) );
  AOI22CDNM1P U100 ( .A(n27), .B(n185), .C(\Queue[4][17] ), .D(n27), .Z(n405)
         );
  AOI22CDNM1P U101 ( .A(n27), .B(n187), .C(\Queue[4][18] ), .D(n27), .Z(n406)
         );
  N1M1P U102 ( .A(Packet_In[19]), .Z(n189) );
  AOI22CDNM1P U103 ( .A(n27), .B(n189), .C(\Queue[4][19] ), .D(n27), .Z(n407)
         );
  AOI22CDNM1P U104 ( .A(n27), .B(n191), .C(\Queue[4][20] ), .D(n27), .Z(n408)
         );
  N1M1P U105 ( .A(Packet_In[21]), .Z(n193) );
  AOI22CDNM1P U106 ( .A(n27), .B(n193), .C(\Queue[4][21] ), .D(n27), .Z(n409)
         );
  AOI22CDNM1P U107 ( .A(n27), .B(n195), .C(\Queue[4][22] ), .D(n27), .Z(n410)
         );
  AOI22CDNM1P U108 ( .A(n27), .B(n197), .C(\Queue[4][23] ), .D(n27), .Z(n411)
         );
  N1M1P U109 ( .A(Packet_In[24]), .Z(n199) );
  AOI22CDNM1P U110 ( .A(n27), .B(n199), .C(\Queue[4][24] ), .D(n27), .Z(n412)
         );
  AOI22CDNM1P U111 ( .A(n27), .B(n201), .C(\Queue[4][25] ), .D(n27), .Z(n413)
         );
  N1M1P U112 ( .A(Packet_In[26]), .Z(n203) );
  AOI22CDNM1P U113 ( .A(n27), .B(n203), .C(\Queue[4][26] ), .D(n27), .Z(n414)
         );
  AOI22CDNM1P U114 ( .A(n27), .B(n205), .C(\Queue[4][27] ), .D(n27), .Z(n415)
         );
  N1M1P U115 ( .A(Packet_In[28]), .Z(n207) );
  AOI22CDNM1P U116 ( .A(n27), .B(n207), .C(\Queue[4][28] ), .D(n27), .Z(n416)
         );
  AOI22CDNM1P U117 ( .A(n27), .B(n373), .C(\Queue[4][29] ), .D(n27), .Z(n417)
         );
  AOI22CDNM1P U118 ( .A(n27), .B(n375), .C(\Queue[4][30] ), .D(n27), .Z(n418)
         );
  OAI22CDNM1P U119 ( .A(n146), .B(n28), .C(n381), .D(Full), .Z(n419) );
  OA21M1P U120 ( .A(n146), .B(n383), .C(n19), .Z(n31) );
  AOI22M1P U121 ( .A(\Queue[2][0] ), .B(n10), .C(\Queue[1][0] ), .D(n7), .Z(
        n32) );
  OAI21M1P U122 ( .A(n151), .B(n66), .C(n32), .Z(n420) );
  AOI22M1P U123 ( .A(n9), .B(\Queue[2][1] ), .C(\Queue[1][1] ), .D(n7), .Z(n33) );
  OAI21M1P U124 ( .A(n66), .B(n153), .C(n33), .Z(n421) );
  AOI22M1P U125 ( .A(n10), .B(\Queue[2][2] ), .C(\Queue[1][2] ), .D(n7), .Z(
        n34) );
  OAI21M1P U126 ( .A(n66), .B(n155), .C(n34), .Z(n422) );
  AOI22M1P U127 ( .A(n10), .B(\Queue[2][3] ), .C(\Queue[1][3] ), .D(n7), .Z(
        n35) );
  OAI21M1P U128 ( .A(n66), .B(n157), .C(n35), .Z(n423) );
  AOI22M1P U129 ( .A(n10), .B(\Queue[2][4] ), .C(\Queue[1][4] ), .D(n7), .Z(
        n36) );
  OAI21M1P U130 ( .A(n66), .B(n159), .C(n36), .Z(n424) );
  AOI22M1P U131 ( .A(n10), .B(\Queue[2][5] ), .C(\Queue[1][5] ), .D(n7), .Z(
        n37) );
  OAI21M1P U132 ( .A(n66), .B(n161), .C(n37), .Z(n425) );
  AOI22M1P U133 ( .A(n10), .B(\Queue[2][6] ), .C(\Queue[1][6] ), .D(n7), .Z(
        n38) );
  OAI21M1P U134 ( .A(n66), .B(n163), .C(n38), .Z(n426) );
  AOI22M1P U135 ( .A(n10), .B(\Queue[2][7] ), .C(\Queue[1][7] ), .D(n7), .Z(
        n39) );
  OAI21M1P U136 ( .A(n66), .B(n165), .C(n39), .Z(n427) );
  AOI22M1P U137 ( .A(n10), .B(\Queue[2][8] ), .C(\Queue[1][8] ), .D(n7), .Z(
        n40) );
  OAI21M1P U138 ( .A(n66), .B(n167), .C(n40), .Z(n428) );
  AOI22M1P U139 ( .A(n10), .B(\Queue[2][9] ), .C(\Queue[1][9] ), .D(n63), .Z(
        n41) );
  OAI21M1P U140 ( .A(n66), .B(n169), .C(n41), .Z(n429) );
  AOI22M1P U141 ( .A(n10), .B(\Queue[2][10] ), .C(\Queue[1][10] ), .D(n8), .Z(
        n42) );
  OAI21M1P U142 ( .A(n66), .B(n171), .C(n42), .Z(n430) );
  AOI22M1P U143 ( .A(n10), .B(\Queue[2][11] ), .C(\Queue[1][11] ), .D(n7), .Z(
        n43) );
  OAI21M1P U144 ( .A(n66), .B(n173), .C(n43), .Z(n431) );
  AOI22M1P U145 ( .A(n9), .B(\Queue[2][12] ), .C(\Queue[1][12] ), .D(n63), .Z(
        n44) );
  OAI21M1P U146 ( .A(n66), .B(n175), .C(n44), .Z(n432) );
  AOI22M1P U147 ( .A(n9), .B(\Queue[2][13] ), .C(\Queue[1][13] ), .D(n63), .Z(
        n45) );
  OAI21M1P U148 ( .A(n66), .B(n177), .C(n45), .Z(n433) );
  AOI22M1P U149 ( .A(n9), .B(\Queue[2][14] ), .C(\Queue[1][14] ), .D(n63), .Z(
        n46) );
  OAI21M1P U150 ( .A(n66), .B(n179), .C(n46), .Z(n434) );
  AOI22M1P U151 ( .A(n9), .B(\Queue[2][15] ), .C(\Queue[1][15] ), .D(n63), .Z(
        n47) );
  OAI21M1P U152 ( .A(n66), .B(n181), .C(n47), .Z(n435) );
  AOI22M1P U153 ( .A(n9), .B(\Queue[2][16] ), .C(\Queue[1][16] ), .D(n63), .Z(
        n48) );
  OAI21M1P U154 ( .A(n66), .B(n183), .C(n48), .Z(n436) );
  AOI22M1P U155 ( .A(n9), .B(\Queue[2][17] ), .C(\Queue[1][17] ), .D(n63), .Z(
        n49) );
  OAI21M1P U156 ( .A(n66), .B(n185), .C(n49), .Z(n437) );
  AOI22M1P U157 ( .A(n9), .B(\Queue[2][18] ), .C(\Queue[1][18] ), .D(n8), .Z(
        n50) );
  OAI21M1P U158 ( .A(n66), .B(n187), .C(n50), .Z(n438) );
  AOI22M1P U159 ( .A(n9), .B(\Queue[2][19] ), .C(\Queue[1][19] ), .D(n8), .Z(
        n51) );
  OAI21M1P U160 ( .A(n66), .B(n189), .C(n51), .Z(n439) );
  AOI22M1P U161 ( .A(n9), .B(\Queue[2][20] ), .C(\Queue[1][20] ), .D(n8), .Z(
        n52) );
  OAI21M1P U162 ( .A(n66), .B(n191), .C(n52), .Z(n440) );
  AOI22M1P U163 ( .A(n9), .B(\Queue[2][21] ), .C(\Queue[1][21] ), .D(n8), .Z(
        n53) );
  OAI21M1P U164 ( .A(n66), .B(n193), .C(n53), .Z(n441) );
  AOI22M1P U165 ( .A(n10), .B(\Queue[2][22] ), .C(\Queue[1][22] ), .D(n8), .Z(
        n54) );
  OAI21M1P U166 ( .A(n66), .B(n195), .C(n54), .Z(n442) );
  AOI22M1P U167 ( .A(n9), .B(\Queue[2][23] ), .C(\Queue[1][23] ), .D(n8), .Z(
        n55) );
  OAI21M1P U168 ( .A(n66), .B(n197), .C(n55), .Z(n443) );
  AOI22M1P U169 ( .A(n10), .B(\Queue[2][24] ), .C(\Queue[1][24] ), .D(n8), .Z(
        n56) );
  OAI21M1P U170 ( .A(n66), .B(n199), .C(n56), .Z(n444) );
  AOI22M1P U171 ( .A(n64), .B(\Queue[2][25] ), .C(\Queue[1][25] ), .D(n8), .Z(
        n57) );
  OAI21M1P U172 ( .A(n66), .B(n201), .C(n57), .Z(n445) );
  AOI22M1P U173 ( .A(n64), .B(\Queue[2][26] ), .C(\Queue[1][26] ), .D(n8), .Z(
        n58) );
  OAI21M1P U174 ( .A(n66), .B(n203), .C(n58), .Z(n446) );
  AOI22M1P U175 ( .A(n64), .B(\Queue[2][27] ), .C(\Queue[1][27] ), .D(n8), .Z(
        n59) );
  OAI21M1P U176 ( .A(n66), .B(n205), .C(n59), .Z(n447) );
  AOI22M1P U177 ( .A(n64), .B(\Queue[2][28] ), .C(\Queue[1][28] ), .D(n7), .Z(
        n60) );
  OAI21M1P U178 ( .A(n66), .B(n207), .C(n60), .Z(n448) );
  AOI22M1P U179 ( .A(n64), .B(\Queue[2][29] ), .C(\Queue[1][29] ), .D(n7), .Z(
        n61) );
  OAI21M1P U180 ( .A(n66), .B(n373), .C(n61), .Z(n449) );
  AOI22M1P U181 ( .A(n64), .B(\Queue[2][30] ), .C(\Queue[1][30] ), .D(n8), .Z(
        n62) );
  OAI21M1P U182 ( .A(n66), .B(n375), .C(n62), .Z(n450) );
  AOI22M1P U183 ( .A(n64), .B(\Queue[2][31] ), .C(\Queue[1][31] ), .D(n8), .Z(
        n65) );
  OAI21M1P U184 ( .A(n66), .B(n380), .C(n65), .Z(n451) );
  OAI21M1P U185 ( .A(n68), .B(n67), .C(n148), .Z(n69) );
  AOI21M1P U186 ( .A(n6), .B(n383), .C(n148), .Z(n102) );
  AOI22M1P U187 ( .A(\Queue[1][0] ), .B(n5), .C(n101), .D(Packet_Out[0]), .Z(
        n70) );
  OAI21M1P U188 ( .A(n151), .B(n14), .C(n70), .Z(n452) );
  AOI22M1P U189 ( .A(\Queue[1][1] ), .B(n5), .C(n101), .D(Packet_Out[1]), .Z(
        n71) );
  OAI21M1P U190 ( .A(n153), .B(n104), .C(n71), .Z(n453) );
  AOI22M1P U191 ( .A(\Queue[1][2] ), .B(n5), .C(n101), .D(Packet_Out[2]), .Z(
        n72) );
  OAI21M1P U192 ( .A(n155), .B(n104), .C(n72), .Z(n454) );
  AOI22M1P U193 ( .A(\Queue[1][3] ), .B(n5), .C(n101), .D(Packet_Out[3]), .Z(
        n73) );
  OAI21M1P U194 ( .A(n157), .B(n104), .C(n73), .Z(n455) );
  AOI22M1P U195 ( .A(\Queue[1][4] ), .B(n5), .C(n101), .D(Packet_Out[4]), .Z(
        n74) );
  OAI21M1P U196 ( .A(n159), .B(n104), .C(n74), .Z(n456) );
  AOI22M1P U197 ( .A(\Queue[1][5] ), .B(n5), .C(n101), .D(Packet_Out[5]), .Z(
        n75) );
  OAI21M1P U198 ( .A(n161), .B(n104), .C(n75), .Z(n457) );
  AOI22M1P U199 ( .A(\Queue[1][6] ), .B(n5), .C(n101), .D(Packet_Out[6]), .Z(
        n76) );
  OAI21M1P U200 ( .A(n163), .B(n104), .C(n76), .Z(n458) );
  AOI22M1P U201 ( .A(\Queue[1][7] ), .B(n5), .C(n101), .D(Packet_Out[7]), .Z(
        n77) );
  OAI21M1P U202 ( .A(n165), .B(n13), .C(n77), .Z(n459) );
  AOI22M1P U203 ( .A(\Queue[1][8] ), .B(n5), .C(n101), .D(Packet_Out[8]), .Z(
        n78) );
  OAI21M1P U204 ( .A(n167), .B(n14), .C(n78), .Z(n460) );
  AOI22M1P U205 ( .A(\Queue[1][9] ), .B(n5), .C(n101), .D(Packet_Out[9]), .Z(
        n79) );
  OAI21M1P U206 ( .A(n169), .B(n13), .C(n79), .Z(n461) );
  AOI22M1P U207 ( .A(\Queue[1][10] ), .B(n5), .C(n11), .D(Packet_Out[10]), .Z(
        n80) );
  OAI21M1P U208 ( .A(n171), .B(n13), .C(n80), .Z(n462) );
  AOI22M1P U209 ( .A(\Queue[1][11] ), .B(n5), .C(n11), .D(Packet_Out[11]), .Z(
        n81) );
  OAI21M1P U210 ( .A(n173), .B(n13), .C(n81), .Z(n463) );
  AOI22M1P U211 ( .A(\Queue[1][12] ), .B(n5), .C(n11), .D(Packet_Out[12]), .Z(
        n82) );
  OAI21M1P U212 ( .A(n175), .B(n13), .C(n82), .Z(n464) );
  AOI22M1P U213 ( .A(\Queue[1][13] ), .B(n5), .C(n11), .D(Packet_Out[13]), .Z(
        n83) );
  OAI21M1P U214 ( .A(n177), .B(n13), .C(n83), .Z(n465) );
  AOI22M1P U215 ( .A(\Queue[1][14] ), .B(n5), .C(n11), .D(Packet_Out[14]), .Z(
        n84) );
  OAI21M1P U216 ( .A(n179), .B(n13), .C(n84), .Z(n466) );
  AOI22M1P U217 ( .A(\Queue[1][15] ), .B(n5), .C(n11), .D(Packet_Out[15]), .Z(
        n85) );
  OAI21M1P U218 ( .A(n181), .B(n13), .C(n85), .Z(n467) );
  AOI22M1P U219 ( .A(\Queue[1][16] ), .B(n5), .C(n11), .D(Packet_Out[16]), .Z(
        n86) );
  OAI21M1P U220 ( .A(n183), .B(n13), .C(n86), .Z(n468) );
  AOI22M1P U221 ( .A(\Queue[1][17] ), .B(n5), .C(n11), .D(Packet_Out[17]), .Z(
        n87) );
  OAI21M1P U222 ( .A(n185), .B(n13), .C(n87), .Z(n469) );
  AOI22M1P U223 ( .A(\Queue[1][18] ), .B(n5), .C(n11), .D(Packet_Out[18]), .Z(
        n88) );
  OAI21M1P U224 ( .A(n187), .B(n13), .C(n88), .Z(n470) );
  AOI22M1P U225 ( .A(\Queue[1][19] ), .B(n5), .C(n11), .D(Packet_Out[19]), .Z(
        n89) );
  OAI21M1P U226 ( .A(n189), .B(n13), .C(n89), .Z(n471) );
  AOI22M1P U227 ( .A(\Queue[1][20] ), .B(n5), .C(n12), .D(Packet_Out[20]), .Z(
        n90) );
  OAI21M1P U228 ( .A(n191), .B(n14), .C(n90), .Z(n472) );
  AOI22M1P U229 ( .A(\Queue[1][21] ), .B(n5), .C(n12), .D(Packet_Out[21]), .Z(
        n91) );
  OAI21M1P U230 ( .A(n193), .B(n14), .C(n91), .Z(n473) );
  AOI22M1P U231 ( .A(\Queue[1][22] ), .B(n5), .C(n12), .D(Packet_Out[22]), .Z(
        n92) );
  OAI21M1P U232 ( .A(n195), .B(n14), .C(n92), .Z(n474) );
  AOI22M1P U233 ( .A(\Queue[1][23] ), .B(n5), .C(n12), .D(Packet_Out[23]), .Z(
        n93) );
  OAI21M1P U234 ( .A(n197), .B(n14), .C(n93), .Z(n475) );
  AOI22M1P U235 ( .A(\Queue[1][24] ), .B(n5), .C(n12), .D(Packet_Out[24]), .Z(
        n94) );
  OAI21M1P U236 ( .A(n199), .B(n14), .C(n94), .Z(n476) );
  AOI22M1P U237 ( .A(\Queue[1][25] ), .B(n5), .C(n12), .D(Packet_Out[25]), .Z(
        n95) );
  OAI21M1P U238 ( .A(n201), .B(n14), .C(n95), .Z(n477) );
  AOI22M1P U239 ( .A(\Queue[1][26] ), .B(n5), .C(n12), .D(Packet_Out[26]), .Z(
        n96) );
  OAI21M1P U240 ( .A(n203), .B(n14), .C(n96), .Z(n478) );
  AOI22M1P U241 ( .A(\Queue[1][27] ), .B(n5), .C(n12), .D(Packet_Out[27]), .Z(
        n97) );
  OAI21M1P U242 ( .A(n205), .B(n14), .C(n97), .Z(n479) );
  AOI22M1P U243 ( .A(\Queue[1][28] ), .B(n5), .C(n12), .D(Packet_Out[28]), .Z(
        n98) );
  OAI21M1P U244 ( .A(n207), .B(n14), .C(n98), .Z(n480) );
  AOI22M1P U245 ( .A(\Queue[1][29] ), .B(n5), .C(n12), .D(Packet_Out[29]), .Z(
        n99) );
  OAI21M1P U246 ( .A(n373), .B(n14), .C(n99), .Z(n481) );
  AOI22M1P U247 ( .A(\Queue[1][30] ), .B(n102), .C(n11), .D(Packet_Out[30]), 
        .Z(n100) );
  OAI21M1P U248 ( .A(n375), .B(n13), .C(n100), .Z(n482) );
  AOI22M1P U249 ( .A(\Queue[1][31] ), .B(n102), .C(n12), .D(Packet_Out[31]), 
        .Z(n103) );
  OAI21M1P U250 ( .A(n380), .B(n14), .C(n103), .Z(n483) );
  OA21M1P U251 ( .A(n146), .B(n107), .C(n19), .Z(n105) );
  ND2M1P U252 ( .A(n106), .B(n144), .Z(n145) );
  AOI21M1P U253 ( .A(n6), .B(n147), .C(n148), .Z(n139) );
  AOI22M1P U254 ( .A(\Queue[2][0] ), .B(n140), .C(\Queue[3][0] ), .D(n4), .Z(
        n108) );
  OAI21M1P U255 ( .A(n151), .B(n16), .C(n108), .Z(n484) );
  AOI22M1P U256 ( .A(\Queue[2][1] ), .B(n140), .C(n4), .D(\Queue[3][1] ), .Z(
        n109) );
  OAI21M1P U257 ( .A(n153), .B(n142), .C(n109), .Z(n485) );
  AOI22M1P U258 ( .A(\Queue[2][2] ), .B(n140), .C(n4), .D(\Queue[3][2] ), .Z(
        n110) );
  OAI21M1P U259 ( .A(n155), .B(n142), .C(n110), .Z(n486) );
  AOI22M1P U260 ( .A(\Queue[2][3] ), .B(n140), .C(n4), .D(\Queue[3][3] ), .Z(
        n111) );
  OAI21M1P U261 ( .A(n157), .B(n142), .C(n111), .Z(n487) );
  AOI22M1P U262 ( .A(\Queue[2][4] ), .B(n140), .C(n4), .D(\Queue[3][4] ), .Z(
        n112) );
  OAI21M1P U263 ( .A(n159), .B(n142), .C(n112), .Z(n488) );
  AOI22M1P U264 ( .A(\Queue[2][5] ), .B(n140), .C(n4), .D(\Queue[3][5] ), .Z(
        n113) );
  OAI21M1P U265 ( .A(n161), .B(n142), .C(n113), .Z(n489) );
  AOI22M1P U266 ( .A(\Queue[2][6] ), .B(n140), .C(n4), .D(\Queue[3][6] ), .Z(
        n114) );
  OAI21M1P U267 ( .A(n163), .B(n142), .C(n114), .Z(n490) );
  AOI22M1P U268 ( .A(\Queue[2][7] ), .B(n140), .C(n4), .D(\Queue[3][7] ), .Z(
        n115) );
  OAI21M1P U269 ( .A(n165), .B(n15), .C(n115), .Z(n491) );
  AOI22M1P U270 ( .A(\Queue[2][8] ), .B(n140), .C(n4), .D(\Queue[3][8] ), .Z(
        n116) );
  OAI21M1P U271 ( .A(n167), .B(n16), .C(n116), .Z(n492) );
  AOI22M1P U272 ( .A(\Queue[2][9] ), .B(n140), .C(n4), .D(\Queue[3][9] ), .Z(
        n117) );
  OAI21M1P U273 ( .A(n169), .B(n15), .C(n117), .Z(n493) );
  AOI22M1P U274 ( .A(\Queue[2][10] ), .B(n140), .C(n4), .D(\Queue[3][10] ), 
        .Z(n118) );
  OAI21M1P U275 ( .A(n171), .B(n15), .C(n118), .Z(n494) );
  AOI22M1P U276 ( .A(\Queue[2][11] ), .B(n140), .C(n4), .D(\Queue[3][11] ), 
        .Z(n119) );
  OAI21M1P U277 ( .A(n173), .B(n15), .C(n119), .Z(n495) );
  AOI22M1P U278 ( .A(\Queue[2][12] ), .B(n140), .C(n4), .D(\Queue[3][12] ), 
        .Z(n120) );
  OAI21M1P U279 ( .A(n175), .B(n15), .C(n120), .Z(n496) );
  AOI22M1P U280 ( .A(\Queue[2][13] ), .B(n140), .C(n4), .D(\Queue[3][13] ), 
        .Z(n121) );
  OAI21M1P U281 ( .A(n177), .B(n15), .C(n121), .Z(n497) );
  AOI22M1P U282 ( .A(\Queue[2][14] ), .B(n140), .C(n4), .D(\Queue[3][14] ), 
        .Z(n122) );
  OAI21M1P U283 ( .A(n179), .B(n15), .C(n122), .Z(n498) );
  AOI22M1P U284 ( .A(\Queue[2][15] ), .B(n140), .C(n4), .D(\Queue[3][15] ), 
        .Z(n123) );
  OAI21M1P U285 ( .A(n181), .B(n15), .C(n123), .Z(n499) );
  AOI22M1P U286 ( .A(\Queue[2][16] ), .B(n140), .C(n4), .D(\Queue[3][16] ), 
        .Z(n124) );
  OAI21M1P U287 ( .A(n183), .B(n15), .C(n124), .Z(n500) );
  AOI22M1P U288 ( .A(\Queue[2][17] ), .B(n140), .C(n4), .D(\Queue[3][17] ), 
        .Z(n125) );
  OAI21M1P U289 ( .A(n185), .B(n15), .C(n125), .Z(n501) );
  AOI22M1P U290 ( .A(\Queue[2][18] ), .B(n140), .C(n4), .D(\Queue[3][18] ), 
        .Z(n126) );
  OAI21M1P U291 ( .A(n187), .B(n15), .C(n126), .Z(n502) );
  AOI22M1P U292 ( .A(\Queue[2][19] ), .B(n140), .C(n4), .D(\Queue[3][19] ), 
        .Z(n127) );
  OAI21M1P U293 ( .A(n189), .B(n15), .C(n127), .Z(n503) );
  AOI22M1P U294 ( .A(\Queue[2][20] ), .B(n140), .C(n4), .D(\Queue[3][20] ), 
        .Z(n128) );
  OAI21M1P U295 ( .A(n191), .B(n16), .C(n128), .Z(n504) );
  AOI22M1P U296 ( .A(\Queue[2][21] ), .B(n140), .C(n4), .D(\Queue[3][21] ), 
        .Z(n129) );
  OAI21M1P U297 ( .A(n193), .B(n16), .C(n129), .Z(n505) );
  AOI22M1P U298 ( .A(\Queue[2][22] ), .B(n140), .C(n4), .D(\Queue[3][22] ), 
        .Z(n130) );
  OAI21M1P U299 ( .A(n195), .B(n16), .C(n130), .Z(n506) );
  AOI22M1P U300 ( .A(\Queue[2][23] ), .B(n140), .C(n4), .D(\Queue[3][23] ), 
        .Z(n131) );
  OAI21M1P U301 ( .A(n197), .B(n16), .C(n131), .Z(n507) );
  AOI22M1P U302 ( .A(\Queue[2][24] ), .B(n140), .C(n4), .D(\Queue[3][24] ), 
        .Z(n132) );
  OAI21M1P U303 ( .A(n199), .B(n16), .C(n132), .Z(n508) );
  AOI22M1P U304 ( .A(\Queue[2][25] ), .B(n140), .C(n4), .D(\Queue[3][25] ), 
        .Z(n133) );
  OAI21M1P U305 ( .A(n201), .B(n16), .C(n133), .Z(n509) );
  AOI22M1P U306 ( .A(\Queue[2][26] ), .B(n140), .C(n4), .D(\Queue[3][26] ), 
        .Z(n134) );
  OAI21M1P U307 ( .A(n203), .B(n16), .C(n134), .Z(n510) );
  AOI22M1P U308 ( .A(\Queue[2][27] ), .B(n140), .C(n4), .D(\Queue[3][27] ), 
        .Z(n135) );
  OAI21M1P U309 ( .A(n205), .B(n16), .C(n135), .Z(n511) );
  AOI22M1P U310 ( .A(\Queue[2][28] ), .B(n140), .C(n4), .D(\Queue[3][28] ), 
        .Z(n136) );
  OAI21M1P U311 ( .A(n207), .B(n16), .C(n136), .Z(n512) );
  AOI22M1P U312 ( .A(\Queue[2][29] ), .B(n140), .C(n4), .D(\Queue[3][29] ), 
        .Z(n137) );
  OAI21M1P U313 ( .A(n373), .B(n16), .C(n137), .Z(n513) );
  AOI22M1P U314 ( .A(\Queue[2][30] ), .B(n140), .C(n4), .D(\Queue[3][30] ), 
        .Z(n138) );
  OAI21M1P U315 ( .A(n375), .B(n15), .C(n138), .Z(n514) );
  AOI22M1P U316 ( .A(\Queue[2][31] ), .B(n140), .C(n4), .D(\Queue[3][31] ), 
        .Z(n141) );
  OAI21M1P U317 ( .A(n380), .B(n16), .C(n141), .Z(n515) );
  OA21M1P U318 ( .A(n146), .B(n147), .C(n19), .Z(n143) );
  AOI21M1P U319 ( .A(n6), .B(n149), .C(n148), .Z(n376) );
  AOI22M1P U320 ( .A(\Queue[3][0] ), .B(n377), .C(n3), .D(\Queue[4][0] ), .Z(
        n150) );
  OAI21M1P U321 ( .A(n151), .B(n18), .C(n150), .Z(n516) );
  AOI22M1P U322 ( .A(\Queue[3][1] ), .B(n377), .C(n3), .D(\Queue[4][1] ), .Z(
        n152) );
  OAI21M1P U323 ( .A(n153), .B(n379), .C(n152), .Z(n517) );
  AOI22M1P U324 ( .A(\Queue[3][2] ), .B(n377), .C(n3), .D(\Queue[4][2] ), .Z(
        n154) );
  OAI21M1P U325 ( .A(n155), .B(n379), .C(n154), .Z(n518) );
  AOI22M1P U326 ( .A(\Queue[3][3] ), .B(n377), .C(n3), .D(\Queue[4][3] ), .Z(
        n156) );
  OAI21M1P U327 ( .A(n157), .B(n379), .C(n156), .Z(n519) );
  AOI22M1P U328 ( .A(\Queue[3][4] ), .B(n377), .C(n3), .D(\Queue[4][4] ), .Z(
        n158) );
  OAI21M1P U329 ( .A(n159), .B(n379), .C(n158), .Z(n520) );
  AOI22M1P U330 ( .A(\Queue[3][5] ), .B(n377), .C(n3), .D(\Queue[4][5] ), .Z(
        n160) );
  OAI21M1P U331 ( .A(n161), .B(n379), .C(n160), .Z(n521) );
  AOI22M1P U332 ( .A(\Queue[3][6] ), .B(n377), .C(n3), .D(\Queue[4][6] ), .Z(
        n162) );
  OAI21M1P U333 ( .A(n163), .B(n379), .C(n162), .Z(n522) );
  AOI22M1P U334 ( .A(\Queue[3][7] ), .B(n377), .C(n3), .D(\Queue[4][7] ), .Z(
        n164) );
  OAI21M1P U335 ( .A(n165), .B(n17), .C(n164), .Z(n523) );
  AOI22M1P U336 ( .A(\Queue[3][8] ), .B(n377), .C(n3), .D(\Queue[4][8] ), .Z(
        n166) );
  OAI21M1P U337 ( .A(n167), .B(n18), .C(n166), .Z(n524) );
  AOI22M1P U338 ( .A(\Queue[3][9] ), .B(n377), .C(n3), .D(\Queue[4][9] ), .Z(
        n168) );
  OAI21M1P U339 ( .A(n169), .B(n17), .C(n168), .Z(n525) );
  AOI22M1P U340 ( .A(\Queue[3][10] ), .B(n377), .C(n3), .D(\Queue[4][10] ), 
        .Z(n170) );
  OAI21M1P U341 ( .A(n171), .B(n17), .C(n170), .Z(n526) );
  AOI22M1P U342 ( .A(\Queue[3][11] ), .B(n377), .C(n3), .D(\Queue[4][11] ), 
        .Z(n172) );
  OAI21M1P U343 ( .A(n173), .B(n17), .C(n172), .Z(n527) );
  AOI22M1P U344 ( .A(\Queue[3][12] ), .B(n377), .C(n3), .D(\Queue[4][12] ), 
        .Z(n174) );
  OAI21M1P U345 ( .A(n175), .B(n17), .C(n174), .Z(n528) );
  AOI22M1P U346 ( .A(\Queue[3][13] ), .B(n377), .C(n3), .D(\Queue[4][13] ), 
        .Z(n176) );
  OAI21M1P U347 ( .A(n177), .B(n17), .C(n176), .Z(n529) );
  AOI22M1P U348 ( .A(\Queue[3][14] ), .B(n377), .C(n3), .D(\Queue[4][14] ), 
        .Z(n178) );
  OAI21M1P U349 ( .A(n179), .B(n17), .C(n178), .Z(n530) );
  AOI22M1P U350 ( .A(\Queue[3][15] ), .B(n377), .C(n3), .D(\Queue[4][15] ), 
        .Z(n180) );
  OAI21M1P U351 ( .A(n181), .B(n17), .C(n180), .Z(n531) );
  AOI22M1P U352 ( .A(\Queue[3][16] ), .B(n377), .C(n3), .D(\Queue[4][16] ), 
        .Z(n182) );
  OAI21M1P U353 ( .A(n183), .B(n17), .C(n182), .Z(n532) );
  AOI22M1P U354 ( .A(\Queue[3][17] ), .B(n377), .C(n3), .D(\Queue[4][17] ), 
        .Z(n184) );
  OAI21M1P U355 ( .A(n185), .B(n17), .C(n184), .Z(n533) );
  AOI22M1P U356 ( .A(\Queue[3][18] ), .B(n377), .C(n3), .D(\Queue[4][18] ), 
        .Z(n186) );
  OAI21M1P U357 ( .A(n187), .B(n17), .C(n186), .Z(n534) );
  AOI22M1P U358 ( .A(\Queue[3][19] ), .B(n377), .C(n3), .D(\Queue[4][19] ), 
        .Z(n188) );
  OAI21M1P U359 ( .A(n189), .B(n17), .C(n188), .Z(n535) );
  AOI22M1P U360 ( .A(\Queue[3][20] ), .B(n377), .C(n3), .D(\Queue[4][20] ), 
        .Z(n190) );
  OAI21M1P U361 ( .A(n191), .B(n18), .C(n190), .Z(n536) );
  AOI22M1P U362 ( .A(\Queue[3][21] ), .B(n377), .C(n3), .D(\Queue[4][21] ), 
        .Z(n192) );
  OAI21M1P U363 ( .A(n193), .B(n18), .C(n192), .Z(n537) );
  AOI22M1P U364 ( .A(\Queue[3][22] ), .B(n377), .C(n3), .D(\Queue[4][22] ), 
        .Z(n194) );
  OAI21M1P U365 ( .A(n195), .B(n18), .C(n194), .Z(n538) );
  AOI22M1P U366 ( .A(\Queue[3][23] ), .B(n377), .C(n3), .D(\Queue[4][23] ), 
        .Z(n196) );
  OAI21M1P U367 ( .A(n197), .B(n18), .C(n196), .Z(n539) );
  AOI22M1P U368 ( .A(\Queue[3][24] ), .B(n377), .C(n3), .D(\Queue[4][24] ), 
        .Z(n198) );
  OAI21M1P U369 ( .A(n199), .B(n18), .C(n198), .Z(n540) );
  AOI22M1P U370 ( .A(\Queue[3][25] ), .B(n377), .C(n3), .D(\Queue[4][25] ), 
        .Z(n200) );
  OAI21M1P U371 ( .A(n201), .B(n18), .C(n200), .Z(n541) );
  AOI22M1P U372 ( .A(\Queue[3][26] ), .B(n377), .C(n3), .D(\Queue[4][26] ), 
        .Z(n202) );
  OAI21M1P U373 ( .A(n203), .B(n18), .C(n202), .Z(n542) );
  AOI22M1P U374 ( .A(\Queue[3][27] ), .B(n377), .C(n3), .D(\Queue[4][27] ), 
        .Z(n204) );
  OAI21M1P U375 ( .A(n205), .B(n18), .C(n204), .Z(n543) );
  AOI22M1P U376 ( .A(\Queue[3][28] ), .B(n377), .C(n3), .D(\Queue[4][28] ), 
        .Z(n206) );
  OAI21M1P U377 ( .A(n207), .B(n18), .C(n206), .Z(n544) );
  AOI22M1P U378 ( .A(\Queue[3][29] ), .B(n377), .C(n3), .D(\Queue[4][29] ), 
        .Z(n208) );
  OAI21M1P U379 ( .A(n373), .B(n18), .C(n208), .Z(n545) );
  AOI22M1P U380 ( .A(\Queue[3][30] ), .B(n377), .C(n3), .D(\Queue[4][30] ), 
        .Z(n374) );
  OAI21M1P U381 ( .A(n375), .B(n17), .C(n374), .Z(n546) );
  AOI22M1P U382 ( .A(\Queue[3][31] ), .B(n377), .C(n3), .D(\Queue[4][31] ), 
        .Z(n378) );
  OAI21M1P U383 ( .A(n380), .B(n18), .C(n378), .Z(n547) );
  N1M1P U384 ( .A(n548), .Z(Empty) );
  AOI22M1P U385 ( .A(n383), .B(n382), .C(n381), .D(Empty), .Z(n549) );
endmodule


module Packet_Queue_2 ( Clk_r, Rst_n, Packet_In, Read_Ack, Write_Ack, 
        Packet_Out, Empty, Full );
  input [31:0] Packet_In;
  output [31:0] Packet_Out;
  input Clk_r, Rst_n, Read_Ack, Write_Ack;
  output Empty, Full;
  wire   \Queue[4][31] , \Queue[4][30] , \Queue[4][29] , \Queue[4][28] ,
         \Queue[4][27] , \Queue[4][26] , \Queue[4][25] , \Queue[4][24] ,
         \Queue[4][15] , \Queue[4][14] , \Queue[4][13] , \Queue[4][12] ,
         \Queue[4][11] , \Queue[4][10] , \Queue[4][9] , \Queue[4][8] ,
         \Queue[4][7] , \Queue[4][6] , \Queue[4][5] , \Queue[4][4] ,
         \Queue[4][3] , \Queue[4][2] , \Queue[4][1] , \Queue[4][0] ,
         \Queue[3][31] , \Queue[3][30] , \Queue[3][29] , \Queue[3][28] ,
         \Queue[3][27] , \Queue[3][26] , \Queue[3][25] , \Queue[3][24] ,
         \Queue[3][15] , \Queue[3][14] , \Queue[3][13] , \Queue[3][12] ,
         \Queue[3][11] , \Queue[3][10] , \Queue[3][9] , \Queue[3][8] ,
         \Queue[3][7] , \Queue[3][6] , \Queue[3][5] , \Queue[3][4] ,
         \Queue[3][3] , \Queue[3][2] , \Queue[3][1] , \Queue[3][0] ,
         \Queue[2][31] , \Queue[2][30] , \Queue[2][29] , \Queue[2][28] ,
         \Queue[2][27] , \Queue[2][26] , \Queue[2][25] , \Queue[2][24] ,
         \Queue[2][15] , \Queue[2][14] , \Queue[2][13] , \Queue[2][12] ,
         \Queue[2][11] , \Queue[2][10] , \Queue[2][9] , \Queue[2][8] ,
         \Queue[2][7] , \Queue[2][6] , \Queue[2][5] , \Queue[2][4] ,
         \Queue[2][3] , \Queue[2][2] , \Queue[2][1] , \Queue[2][0] ,
         \Queue[1][31] , \Queue[1][30] , \Queue[1][29] , \Queue[1][28] ,
         \Queue[1][27] , \Queue[1][26] , \Queue[1][25] , \Queue[1][24] ,
         \Queue[1][15] , \Queue[1][14] , \Queue[1][13] , \Queue[1][12] ,
         \Queue[1][11] , \Queue[1][10] , \Queue[1][9] , \Queue[1][8] ,
         \Queue[1][7] , \Queue[1][6] , \Queue[1][5] , \Queue[1][4] ,
         \Queue[1][3] , \Queue[1][2] , \Queue[1][1] , \Queue[1][0] , n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n217, n218, n219, n220,
         n221, n222, n223, n224, n249, n250, n251, n252, n253, n254, n255,
         n256, n281, n282, n283, n284, n285, n286, n287, n288, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364;
  wire   [2:0] Count;

  FDN2QM1P \Count_reg[0]  ( .D(n174), .CPN(Clk_r), .CD(Rst_n), .Q(Count[0]) );
  FDN2QM1P \Count_reg[1]  ( .D(n175), .CPN(Clk_r), .CD(Rst_n), .Q(Count[1]) );
  FDN2QM1P \Count_reg[2]  ( .D(n176), .CPN(Clk_r), .CD(Rst_n), .Q(Count[2]) );
  FDN1QM1P \Queue_reg[4][30]  ( .D(n200), .CPN(Clk_r), .Q(\Queue[4][30] ) );
  FDN1QM1P \Queue_reg[3][30]  ( .D(n361), .CPN(Clk_r), .Q(\Queue[3][30] ) );
  FDN1QM1P \Queue_reg[2][30]  ( .D(n337), .CPN(Clk_r), .Q(\Queue[2][30] ) );
  FDN1QM1P \Queue_reg[4][29]  ( .D(n199), .CPN(Clk_r), .Q(\Queue[4][29] ) );
  FDN1QM1P \Queue_reg[3][29]  ( .D(n360), .CPN(Clk_r), .Q(\Queue[3][29] ) );
  FDN1QM1P \Queue_reg[2][29]  ( .D(n336), .CPN(Clk_r), .Q(\Queue[2][29] ) );
  FDN1QM1P \Queue_reg[4][28]  ( .D(n198), .CPN(Clk_r), .Q(\Queue[4][28] ) );
  FDN1QM1P \Queue_reg[3][28]  ( .D(n359), .CPN(Clk_r), .Q(\Queue[3][28] ) );
  FDN1QM1P \Queue_reg[2][28]  ( .D(n335), .CPN(Clk_r), .Q(\Queue[2][28] ) );
  FDN1QM1P \Queue_reg[4][27]  ( .D(n197), .CPN(Clk_r), .Q(\Queue[4][27] ) );
  FDN1QM1P \Queue_reg[3][27]  ( .D(n358), .CPN(Clk_r), .Q(\Queue[3][27] ) );
  FDN1QM1P \Queue_reg[2][27]  ( .D(n334), .CPN(Clk_r), .Q(\Queue[2][27] ) );
  FDN1QM1P \Queue_reg[4][26]  ( .D(n196), .CPN(Clk_r), .Q(\Queue[4][26] ) );
  FDN1QM1P \Queue_reg[3][26]  ( .D(n357), .CPN(Clk_r), .Q(\Queue[3][26] ) );
  FDN1QM1P \Queue_reg[2][26]  ( .D(n333), .CPN(Clk_r), .Q(\Queue[2][26] ) );
  FDN1QM1P \Queue_reg[4][25]  ( .D(n195), .CPN(Clk_r), .Q(\Queue[4][25] ) );
  FDN1QM1P \Queue_reg[3][25]  ( .D(n356), .CPN(Clk_r), .Q(\Queue[3][25] ) );
  FDN1QM1P \Queue_reg[2][25]  ( .D(n332), .CPN(Clk_r), .Q(\Queue[2][25] ) );
  FDN1QM1P \Queue_reg[4][24]  ( .D(n194), .CPN(Clk_r), .Q(\Queue[4][24] ) );
  FDN1QM1P \Queue_reg[3][24]  ( .D(n355), .CPN(Clk_r), .Q(\Queue[3][24] ) );
  FDN1QM1P \Queue_reg[2][24]  ( .D(n331), .CPN(Clk_r), .Q(\Queue[2][24] ) );
  FDN1QM1P \Queue_reg[4][15]  ( .D(n193), .CPN(Clk_r), .Q(\Queue[4][15] ) );
  FDN1QM1P \Queue_reg[3][15]  ( .D(n354), .CPN(Clk_r), .Q(\Queue[3][15] ) );
  FDN1QM1P \Queue_reg[2][15]  ( .D(n330), .CPN(Clk_r), .Q(\Queue[2][15] ) );
  FDN1QM1P \Queue_reg[4][14]  ( .D(n192), .CPN(Clk_r), .Q(\Queue[4][14] ) );
  FDN1QM1P \Queue_reg[3][14]  ( .D(n353), .CPN(Clk_r), .Q(\Queue[3][14] ) );
  FDN1QM1P \Queue_reg[2][14]  ( .D(n329), .CPN(Clk_r), .Q(\Queue[2][14] ) );
  FDN1QM1P \Queue_reg[4][13]  ( .D(n191), .CPN(Clk_r), .Q(\Queue[4][13] ) );
  FDN1QM1P \Queue_reg[3][13]  ( .D(n352), .CPN(Clk_r), .Q(\Queue[3][13] ) );
  FDN1QM1P \Queue_reg[2][13]  ( .D(n328), .CPN(Clk_r), .Q(\Queue[2][13] ) );
  FDN1QM1P \Queue_reg[4][12]  ( .D(n190), .CPN(Clk_r), .Q(\Queue[4][12] ) );
  FDN1QM1P \Queue_reg[3][12]  ( .D(n351), .CPN(Clk_r), .Q(\Queue[3][12] ) );
  FDN1QM1P \Queue_reg[2][12]  ( .D(n327), .CPN(Clk_r), .Q(\Queue[2][12] ) );
  FDN1QM1P \Queue_reg[4][11]  ( .D(n189), .CPN(Clk_r), .Q(\Queue[4][11] ) );
  FDN1QM1P \Queue_reg[3][11]  ( .D(n350), .CPN(Clk_r), .Q(\Queue[3][11] ) );
  FDN1QM1P \Queue_reg[2][11]  ( .D(n326), .CPN(Clk_r), .Q(\Queue[2][11] ) );
  FDN1QM1P \Queue_reg[4][10]  ( .D(n188), .CPN(Clk_r), .Q(\Queue[4][10] ) );
  FDN1QM1P \Queue_reg[3][10]  ( .D(n349), .CPN(Clk_r), .Q(\Queue[3][10] ) );
  FDN1QM1P \Queue_reg[2][10]  ( .D(n325), .CPN(Clk_r), .Q(\Queue[2][10] ) );
  FDN1QM1P \Queue_reg[4][9]  ( .D(n187), .CPN(Clk_r), .Q(\Queue[4][9] ) );
  FDN1QM1P \Queue_reg[3][9]  ( .D(n348), .CPN(Clk_r), .Q(\Queue[3][9] ) );
  FDN1QM1P \Queue_reg[2][9]  ( .D(n324), .CPN(Clk_r), .Q(\Queue[2][9] ) );
  FDN1QM1P \Queue_reg[4][8]  ( .D(n186), .CPN(Clk_r), .Q(\Queue[4][8] ) );
  FDN1QM1P \Queue_reg[3][8]  ( .D(n347), .CPN(Clk_r), .Q(\Queue[3][8] ) );
  FDN1QM1P \Queue_reg[2][8]  ( .D(n323), .CPN(Clk_r), .Q(\Queue[2][8] ) );
  FDN1QM1P \Queue_reg[4][7]  ( .D(n185), .CPN(Clk_r), .Q(\Queue[4][7] ) );
  FDN1QM1P \Queue_reg[3][7]  ( .D(n346), .CPN(Clk_r), .Q(\Queue[3][7] ) );
  FDN1QM1P \Queue_reg[2][7]  ( .D(n322), .CPN(Clk_r), .Q(\Queue[2][7] ) );
  FDN1QM1P \Queue_reg[4][6]  ( .D(n184), .CPN(Clk_r), .Q(\Queue[4][6] ) );
  FDN1QM1P \Queue_reg[3][6]  ( .D(n345), .CPN(Clk_r), .Q(\Queue[3][6] ) );
  FDN1QM1P \Queue_reg[2][6]  ( .D(n321), .CPN(Clk_r), .Q(\Queue[2][6] ) );
  FDN1QM1P \Queue_reg[4][5]  ( .D(n183), .CPN(Clk_r), .Q(\Queue[4][5] ) );
  FDN1QM1P \Queue_reg[3][5]  ( .D(n344), .CPN(Clk_r), .Q(\Queue[3][5] ) );
  FDN1QM1P \Queue_reg[2][5]  ( .D(n320), .CPN(Clk_r), .Q(\Queue[2][5] ) );
  FDN1QM1P \Queue_reg[4][4]  ( .D(n182), .CPN(Clk_r), .Q(\Queue[4][4] ) );
  FDN1QM1P \Queue_reg[3][4]  ( .D(n343), .CPN(Clk_r), .Q(\Queue[3][4] ) );
  FDN1QM1P \Queue_reg[2][4]  ( .D(n319), .CPN(Clk_r), .Q(\Queue[2][4] ) );
  FDN1QM1P \Queue_reg[4][3]  ( .D(n181), .CPN(Clk_r), .Q(\Queue[4][3] ) );
  FDN1QM1P \Queue_reg[3][3]  ( .D(n342), .CPN(Clk_r), .Q(\Queue[3][3] ) );
  FDN1QM1P \Queue_reg[2][3]  ( .D(n318), .CPN(Clk_r), .Q(\Queue[2][3] ) );
  FDN1QM1P \Queue_reg[4][2]  ( .D(n180), .CPN(Clk_r), .Q(\Queue[4][2] ) );
  FDN1QM1P \Queue_reg[3][2]  ( .D(n341), .CPN(Clk_r), .Q(\Queue[3][2] ) );
  FDN1QM1P \Queue_reg[2][2]  ( .D(n317), .CPN(Clk_r), .Q(\Queue[2][2] ) );
  FDN1QM1P \Queue_reg[4][1]  ( .D(n179), .CPN(Clk_r), .Q(\Queue[4][1] ) );
  FDN1QM1P \Queue_reg[3][1]  ( .D(n340), .CPN(Clk_r), .Q(\Queue[3][1] ) );
  FDN1QM1P \Queue_reg[2][1]  ( .D(n316), .CPN(Clk_r), .Q(\Queue[2][1] ) );
  FDN1QM1P \Queue_reg[4][0]  ( .D(n178), .CPN(Clk_r), .Q(\Queue[4][0] ) );
  FDN1QM1P \Queue_reg[3][0]  ( .D(n339), .CPN(Clk_r), .Q(\Queue[3][0] ) );
  FDN1QM1P \Queue_reg[2][0]  ( .D(n315), .CPN(Clk_r), .Q(\Queue[2][0] ) );
  FDN1QM1P \Queue_reg[4][31]  ( .D(n177), .CPN(Clk_r), .Q(\Queue[4][31] ) );
  FDN1QM1P \Queue_reg[3][31]  ( .D(n362), .CPN(Clk_r), .Q(\Queue[3][31] ) );
  FDN1QM1P \Queue_reg[2][31]  ( .D(n338), .CPN(Clk_r), .Q(\Queue[2][31] ) );
  FDN2QM1P Full_reg ( .D(n201), .CPN(Clk_r), .CD(Rst_n), .Q(Full) );
  FDN1QM1P \Queue_reg[1][31]  ( .D(n281), .CPN(Clk_r), .Q(\Queue[1][31] ) );
  FDN1QM1P \Queue_reg[0][31]  ( .D(n314), .CPN(Clk_r), .Q(Packet_Out[31]) );
  FDN1QM1P \Queue_reg[1][30]  ( .D(n256), .CPN(Clk_r), .Q(\Queue[1][30] ) );
  FDN1QM1P \Queue_reg[0][30]  ( .D(n313), .CPN(Clk_r), .Q(Packet_Out[30]) );
  FDN1QM1P \Queue_reg[1][29]  ( .D(n255), .CPN(Clk_r), .Q(\Queue[1][29] ) );
  FDN1QM1P \Queue_reg[0][29]  ( .D(n312), .CPN(Clk_r), .Q(Packet_Out[29]) );
  FDN1QM1P \Queue_reg[1][28]  ( .D(n254), .CPN(Clk_r), .Q(\Queue[1][28] ) );
  FDN1QM1P \Queue_reg[0][28]  ( .D(n311), .CPN(Clk_r), .Q(Packet_Out[28]) );
  FDN1QM1P \Queue_reg[1][27]  ( .D(n253), .CPN(Clk_r), .Q(\Queue[1][27] ) );
  FDN1QM1P \Queue_reg[0][27]  ( .D(n310), .CPN(Clk_r), .Q(Packet_Out[27]) );
  FDN1QM1P \Queue_reg[1][26]  ( .D(n252), .CPN(Clk_r), .Q(\Queue[1][26] ) );
  FDN1QM1P \Queue_reg[0][26]  ( .D(n309), .CPN(Clk_r), .Q(Packet_Out[26]) );
  FDN1QM1P \Queue_reg[1][25]  ( .D(n251), .CPN(Clk_r), .Q(\Queue[1][25] ) );
  FDN1QM1P \Queue_reg[0][25]  ( .D(n308), .CPN(Clk_r), .Q(Packet_Out[25]) );
  FDN1QM1P \Queue_reg[1][24]  ( .D(n250), .CPN(Clk_r), .Q(\Queue[1][24] ) );
  FDN1QM1P \Queue_reg[0][24]  ( .D(n307), .CPN(Clk_r), .Q(Packet_Out[24]) );
  FDN1QM1P \Queue_reg[1][15]  ( .D(n249), .CPN(Clk_r), .Q(\Queue[1][15] ) );
  FDN1QM1P \Queue_reg[0][15]  ( .D(n306), .CPN(Clk_r), .Q(Packet_Out[15]) );
  FDN1QM1P \Queue_reg[1][14]  ( .D(n224), .CPN(Clk_r), .Q(\Queue[1][14] ) );
  FDN1QM1P \Queue_reg[0][14]  ( .D(n305), .CPN(Clk_r), .Q(Packet_Out[14]) );
  FDN1QM1P \Queue_reg[1][13]  ( .D(n223), .CPN(Clk_r), .Q(\Queue[1][13] ) );
  FDN1QM1P \Queue_reg[0][13]  ( .D(n304), .CPN(Clk_r), .Q(Packet_Out[13]) );
  FDN1QM1P \Queue_reg[1][12]  ( .D(n222), .CPN(Clk_r), .Q(\Queue[1][12] ) );
  FDN1QM1P \Queue_reg[0][12]  ( .D(n303), .CPN(Clk_r), .Q(Packet_Out[12]) );
  FDN1QM1P \Queue_reg[1][11]  ( .D(n221), .CPN(Clk_r), .Q(\Queue[1][11] ) );
  FDN1QM1P \Queue_reg[0][11]  ( .D(n302), .CPN(Clk_r), .Q(Packet_Out[11]) );
  FDN1QM1P \Queue_reg[1][10]  ( .D(n220), .CPN(Clk_r), .Q(\Queue[1][10] ) );
  FDN1QM1P \Queue_reg[0][10]  ( .D(n301), .CPN(Clk_r), .Q(Packet_Out[10]) );
  FDN1QM1P \Queue_reg[1][9]  ( .D(n219), .CPN(Clk_r), .Q(\Queue[1][9] ) );
  FDN1QM1P \Queue_reg[0][9]  ( .D(n300), .CPN(Clk_r), .Q(Packet_Out[9]) );
  FDN1QM1P \Queue_reg[1][8]  ( .D(n218), .CPN(Clk_r), .Q(\Queue[1][8] ) );
  FDN1QM1P \Queue_reg[0][8]  ( .D(n299), .CPN(Clk_r), .Q(Packet_Out[8]) );
  FDN1QM1P \Queue_reg[1][7]  ( .D(n217), .CPN(Clk_r), .Q(\Queue[1][7] ) );
  FDN1QM1P \Queue_reg[0][7]  ( .D(n298), .CPN(Clk_r), .Q(Packet_Out[7]) );
  FDN1QM1P \Queue_reg[1][6]  ( .D(n208), .CPN(Clk_r), .Q(\Queue[1][6] ) );
  FDN1QM1P \Queue_reg[0][6]  ( .D(n288), .CPN(Clk_r), .Q(Packet_Out[6]) );
  FDN1QM1P \Queue_reg[1][5]  ( .D(n207), .CPN(Clk_r), .Q(\Queue[1][5] ) );
  FDN1QM1P \Queue_reg[0][5]  ( .D(n287), .CPN(Clk_r), .Q(Packet_Out[5]) );
  FDN1QM1P \Queue_reg[1][4]  ( .D(n206), .CPN(Clk_r), .Q(\Queue[1][4] ) );
  FDN1QM1P \Queue_reg[0][4]  ( .D(n286), .CPN(Clk_r), .Q(Packet_Out[4]) );
  FDN1QM1P \Queue_reg[1][3]  ( .D(n205), .CPN(Clk_r), .Q(\Queue[1][3] ) );
  FDN1QM1P \Queue_reg[0][3]  ( .D(n285), .CPN(Clk_r), .Q(Packet_Out[3]) );
  FDN1QM1P \Queue_reg[1][2]  ( .D(n204), .CPN(Clk_r), .Q(\Queue[1][2] ) );
  FDN1QM1P \Queue_reg[0][2]  ( .D(n284), .CPN(Clk_r), .Q(Packet_Out[2]) );
  FDN1QM1P \Queue_reg[1][1]  ( .D(n203), .CPN(Clk_r), .Q(\Queue[1][1] ) );
  FDN1QM1P \Queue_reg[0][1]  ( .D(n283), .CPN(Clk_r), .Q(Packet_Out[1]) );
  FDN1QM1P \Queue_reg[1][0]  ( .D(n202), .CPN(Clk_r), .Q(\Queue[1][0] ) );
  FDN1QM1P \Queue_reg[0][0]  ( .D(n282), .CPN(Clk_r), .Q(Packet_Out[0]) );
  FDN2QM1P Empty_reg ( .D(n364), .CPN(Clk_r), .CD(Rst_n), .Q(n363) );
  ND2M1P U3 ( .A(Read_Ack), .B(Rst_n), .Z(n118) );
  ND2M1P U4 ( .A(n19), .B(Rst_n), .Z(n54) );
  N1M1P U5 ( .A(n363), .Z(Empty) );
  BUFM2P U6 ( .A(n80), .Z(n11) );
  BUFM2P U7 ( .A(n50), .Z(n8) );
  BUFM2P U8 ( .A(n52), .Z(n5) );
  BUFM2P U9 ( .A(n167), .Z(n13) );
  BUFM2P U10 ( .A(n110), .Z(n7) );
  BUFM2P U11 ( .A(n109), .Z(n9) );
  BUFM2P U12 ( .A(n112), .Z(n3) );
  BUFM2P U13 ( .A(n166), .Z(n10) );
  BUFM2P U14 ( .A(n169), .Z(n4) );
  N1M1P U15 ( .A(Read_Ack), .Z(n114) );
  OAI211M4P U16 ( .A(n173), .B(n114), .C(n12), .D(n55), .Z(n82) );
  N1M2P U17 ( .A(n55), .Z(n79) );
  OAI21M2P U18 ( .A(n12), .B(Read_Ack), .C(n25), .Z(n49) );
  BUFM2P U19 ( .A(n49), .Z(n6) );
  NR3M1P U20 ( .A(Count[0]), .B(Count[1]), .C(n20), .Z(n119) );
  N1M1P U21 ( .A(n119), .Z(n22) );
  NR3M1P U22 ( .A(Count[0]), .B(Count[2]), .C(n23), .Z(n85) );
  NR3M1P U23 ( .A(n24), .B(Count[2]), .C(Count[1]), .Z(n173) );
  NR3M1P U24 ( .A(Count[2]), .B(n24), .C(n23), .Z(n117) );
  N1M1P U25 ( .A(Count[0]), .Z(n24) );
  N1M1P U26 ( .A(Count[2]), .Z(n20) );
  N1M1P U27 ( .A(Count[1]), .Z(n23) );
  NR2FM2P U28 ( .A(n54), .B(n22), .Z(n21) );
  NR2M3P U29 ( .A(Read_Ack), .B(n84), .Z(n19) );
  BUFM3P U30 ( .A(Write_Ack), .Z(n12) );
  N1M1P U31 ( .A(Packet_In[29]), .Z(n163) );
  N1M1P U32 ( .A(Packet_In[28]), .Z(n161) );
  N1M1P U33 ( .A(Packet_In[14]), .Z(n149) );
  N1M1P U34 ( .A(Packet_In[8]), .Z(n137) );
  N1M1P U35 ( .A(Packet_In[10]), .Z(n141) );
  N1M1P U36 ( .A(Packet_In[24]), .Z(n153) );
  N1M1P U37 ( .A(Packet_In[12]), .Z(n145) );
  N1M1P U38 ( .A(Packet_In[15]), .Z(n151) );
  N1M1P U39 ( .A(Packet_In[26]), .Z(n157) );
  N1M1P U40 ( .A(Packet_In[30]), .Z(n165) );
  N1M1P U41 ( .A(Packet_In[4]), .Z(n129) );
  N1M1P U42 ( .A(Packet_In[5]), .Z(n131) );
  N1M1P U43 ( .A(Packet_In[7]), .Z(n135) );
  N1M1P U44 ( .A(Packet_In[2]), .Z(n125) );
  N1M1P U45 ( .A(Packet_In[25]), .Z(n155) );
  N1M1P U46 ( .A(Packet_In[1]), .Z(n123) );
  N1M1P U47 ( .A(Packet_In[13]), .Z(n147) );
  N1M1P U48 ( .A(Packet_In[3]), .Z(n127) );
  N1M1P U49 ( .A(Packet_In[9]), .Z(n139) );
  N1M1P U50 ( .A(Packet_In[31]), .Z(n170) );
  N1M1P U51 ( .A(Packet_In[0]), .Z(n121) );
  N1M1P U52 ( .A(Packet_In[6]), .Z(n133) );
  N1M1P U53 ( .A(Packet_In[27]), .Z(n159) );
  N1M1P U54 ( .A(Packet_In[11]), .Z(n143) );
  N1M2P U55 ( .A(n12), .Z(n84) );
  OAI211M1P U56 ( .A(n85), .B(n116), .C(Rst_n), .D(n115), .Z(n110) );
  OAI211M1P U57 ( .A(n117), .B(n116), .C(Rst_n), .D(n115), .Z(n167) );
  N1M2P U58 ( .A(n19), .Z(n116) );
  NR2M1P U59 ( .A(n114), .B(n12), .Z(n172) );
  NR2M1P U60 ( .A(n19), .B(n172), .Z(n171) );
  AOI22CDNM1P U61 ( .A(n171), .B(n24), .C(n171), .D(n24), .Z(n174) );
  N1M1P U62 ( .A(n172), .Z(n18) );
  AOI22M1P U63 ( .A(Count[0]), .B(n116), .C(n18), .D(n24), .Z(n15) );
  AOI22CDNM1P U64 ( .A(Count[1]), .B(n15), .C(n15), .D(Count[1]), .Z(n175) );
  ND3M1P U65 ( .A(n24), .B(n20), .C(n23), .Z(n53) );
  ND2M1P U66 ( .A(Count[1]), .B(Read_Ack), .Z(n14) );
  OAI211M1P U67 ( .A(Count[1]), .B(n116), .C(n15), .D(n14), .Z(n16) );
  AOI22M1P U68 ( .A(n19), .B(n117), .C(Count[2]), .D(n16), .Z(n17) );
  OAI21M1P U69 ( .A(n53), .B(n18), .C(n17), .Z(n176) );
  AOI22CDNM1P U70 ( .A(n21), .B(n170), .C(\Queue[4][31] ), .D(n21), .Z(n177)
         );
  AOI22CDNM1P U71 ( .A(n21), .B(n121), .C(\Queue[4][0] ), .D(n21), .Z(n178) );
  AOI22CDNM1P U72 ( .A(n21), .B(n123), .C(\Queue[4][1] ), .D(n21), .Z(n179) );
  AOI22CDNM1P U73 ( .A(n21), .B(n125), .C(\Queue[4][2] ), .D(n21), .Z(n180) );
  AOI22CDNM1P U74 ( .A(n21), .B(n127), .C(\Queue[4][3] ), .D(n21), .Z(n181) );
  AOI22CDNM1P U75 ( .A(n21), .B(n129), .C(\Queue[4][4] ), .D(n21), .Z(n182) );
  AOI22CDNM1P U76 ( .A(n21), .B(n131), .C(\Queue[4][5] ), .D(n21), .Z(n183) );
  AOI22CDNM1P U77 ( .A(n21), .B(n133), .C(\Queue[4][6] ), .D(n21), .Z(n184) );
  AOI22CDNM1P U78 ( .A(n21), .B(n135), .C(\Queue[4][7] ), .D(n21), .Z(n185) );
  AOI22CDNM1P U79 ( .A(n21), .B(n137), .C(\Queue[4][8] ), .D(n21), .Z(n186) );
  AOI22CDNM1P U80 ( .A(n21), .B(n139), .C(\Queue[4][9] ), .D(n21), .Z(n187) );
  AOI22CDNM1P U81 ( .A(n21), .B(n141), .C(\Queue[4][10] ), .D(n21), .Z(n188)
         );
  AOI22CDNM1P U82 ( .A(n21), .B(n143), .C(\Queue[4][11] ), .D(n21), .Z(n189)
         );
  AOI22CDNM1P U83 ( .A(n21), .B(n145), .C(\Queue[4][12] ), .D(n21), .Z(n190)
         );
  AOI22CDNM1P U84 ( .A(n21), .B(n147), .C(\Queue[4][13] ), .D(n21), .Z(n191)
         );
  AOI22CDNM1P U85 ( .A(n21), .B(n149), .C(\Queue[4][14] ), .D(n21), .Z(n192)
         );
  AOI22CDNM1P U86 ( .A(n21), .B(n151), .C(\Queue[4][15] ), .D(n21), .Z(n193)
         );
  AOI22CDNM1P U87 ( .A(n21), .B(n153), .C(\Queue[4][24] ), .D(n21), .Z(n194)
         );
  AOI22CDNM1P U88 ( .A(n21), .B(n155), .C(\Queue[4][25] ), .D(n21), .Z(n195)
         );
  AOI22CDNM1P U89 ( .A(n21), .B(n157), .C(\Queue[4][26] ), .D(n21), .Z(n196)
         );
  AOI22CDNM1P U90 ( .A(n21), .B(n159), .C(\Queue[4][27] ), .D(n21), .Z(n197)
         );
  AOI22CDNM1P U91 ( .A(n21), .B(n161), .C(\Queue[4][28] ), .D(n21), .Z(n198)
         );
  AOI22CDNM1P U92 ( .A(n21), .B(n163), .C(\Queue[4][29] ), .D(n21), .Z(n199)
         );
  AOI22CDNM1P U93 ( .A(n21), .B(n165), .C(\Queue[4][30] ), .D(n21), .Z(n200)
         );
  OAI22CDNM1P U94 ( .A(n116), .B(n22), .C(n171), .D(Full), .Z(n201) );
  OA21M1P U95 ( .A(n116), .B(n173), .C(Rst_n), .Z(n25) );
  OAI211M1P U96 ( .A(n85), .B(n114), .C(n12), .D(n25), .Z(n52) );
  AOI21M1P U97 ( .A(n12), .B(n85), .C(n118), .Z(n50) );
  AOI22M1P U98 ( .A(\Queue[2][0] ), .B(n8), .C(\Queue[1][0] ), .D(n6), .Z(n26)
         );
  OAI21M1P U99 ( .A(n121), .B(n5), .C(n26), .Z(n202) );
  AOI22M1P U100 ( .A(n8), .B(\Queue[2][1] ), .C(\Queue[1][1] ), .D(n6), .Z(n27) );
  OAI21M1P U101 ( .A(n5), .B(n123), .C(n27), .Z(n203) );
  AOI22M1P U102 ( .A(n8), .B(\Queue[2][2] ), .C(\Queue[1][2] ), .D(n6), .Z(n28) );
  OAI21M1P U103 ( .A(n5), .B(n125), .C(n28), .Z(n204) );
  AOI22M1P U104 ( .A(n8), .B(\Queue[2][3] ), .C(\Queue[1][3] ), .D(n6), .Z(n29) );
  OAI21M1P U105 ( .A(n5), .B(n127), .C(n29), .Z(n205) );
  AOI22M1P U106 ( .A(n8), .B(\Queue[2][4] ), .C(\Queue[1][4] ), .D(n6), .Z(n30) );
  OAI21M1P U107 ( .A(n5), .B(n129), .C(n30), .Z(n206) );
  AOI22M1P U108 ( .A(n8), .B(\Queue[2][5] ), .C(\Queue[1][5] ), .D(n6), .Z(n31) );
  OAI21M1P U109 ( .A(n5), .B(n131), .C(n31), .Z(n207) );
  AOI22M1P U110 ( .A(n8), .B(\Queue[2][6] ), .C(\Queue[1][6] ), .D(n6), .Z(n32) );
  OAI21M1P U111 ( .A(n5), .B(n133), .C(n32), .Z(n208) );
  AOI22M1P U112 ( .A(n8), .B(\Queue[2][7] ), .C(\Queue[1][7] ), .D(n6), .Z(n33) );
  OAI21M1P U113 ( .A(n5), .B(n135), .C(n33), .Z(n217) );
  AOI22M1P U114 ( .A(n8), .B(\Queue[2][8] ), .C(\Queue[1][8] ), .D(n6), .Z(n34) );
  OAI21M1P U115 ( .A(n5), .B(n137), .C(n34), .Z(n218) );
  AOI22M1P U116 ( .A(n8), .B(\Queue[2][9] ), .C(\Queue[1][9] ), .D(n49), .Z(
        n35) );
  OAI21M1P U117 ( .A(n5), .B(n139), .C(n35), .Z(n219) );
  AOI22M1P U118 ( .A(n8), .B(\Queue[2][10] ), .C(\Queue[1][10] ), .D(n49), .Z(
        n36) );
  OAI21M1P U119 ( .A(n5), .B(n141), .C(n36), .Z(n220) );
  AOI22M1P U120 ( .A(n8), .B(\Queue[2][11] ), .C(\Queue[1][11] ), .D(n49), .Z(
        n37) );
  OAI21M1P U121 ( .A(n5), .B(n143), .C(n37), .Z(n221) );
  AOI22M1P U122 ( .A(n8), .B(\Queue[2][12] ), .C(\Queue[1][12] ), .D(n49), .Z(
        n38) );
  OAI21M1P U123 ( .A(n5), .B(n145), .C(n38), .Z(n222) );
  AOI22M1P U124 ( .A(n8), .B(\Queue[2][13] ), .C(\Queue[1][13] ), .D(n49), .Z(
        n39) );
  OAI21M1P U125 ( .A(n5), .B(n147), .C(n39), .Z(n223) );
  AOI22M1P U126 ( .A(n8), .B(\Queue[2][14] ), .C(\Queue[1][14] ), .D(n49), .Z(
        n40) );
  OAI21M1P U127 ( .A(n5), .B(n149), .C(n40), .Z(n224) );
  AOI22M1P U128 ( .A(n8), .B(\Queue[2][15] ), .C(\Queue[1][15] ), .D(n49), .Z(
        n41) );
  OAI21M1P U129 ( .A(n5), .B(n151), .C(n41), .Z(n249) );
  AOI22M1P U130 ( .A(n8), .B(\Queue[2][24] ), .C(\Queue[1][24] ), .D(n6), .Z(
        n42) );
  OAI21M1P U131 ( .A(n5), .B(n153), .C(n42), .Z(n250) );
  AOI22M1P U132 ( .A(n8), .B(\Queue[2][25] ), .C(\Queue[1][25] ), .D(n6), .Z(
        n43) );
  OAI21M1P U133 ( .A(n5), .B(n155), .C(n43), .Z(n251) );
  AOI22M1P U134 ( .A(n8), .B(\Queue[2][26] ), .C(\Queue[1][26] ), .D(n6), .Z(
        n44) );
  OAI21M1P U135 ( .A(n5), .B(n157), .C(n44), .Z(n252) );
  AOI22M1P U136 ( .A(n8), .B(\Queue[2][27] ), .C(\Queue[1][27] ), .D(n6), .Z(
        n45) );
  OAI21M1P U137 ( .A(n5), .B(n159), .C(n45), .Z(n253) );
  AOI22M1P U138 ( .A(n8), .B(\Queue[2][28] ), .C(\Queue[1][28] ), .D(n6), .Z(
        n46) );
  OAI21M1P U139 ( .A(n5), .B(n161), .C(n46), .Z(n254) );
  AOI22M1P U140 ( .A(n8), .B(\Queue[2][29] ), .C(\Queue[1][29] ), .D(n6), .Z(
        n47) );
  OAI21M1P U141 ( .A(n5), .B(n163), .C(n47), .Z(n255) );
  AOI22M1P U142 ( .A(n8), .B(\Queue[2][30] ), .C(\Queue[1][30] ), .D(n6), .Z(
        n48) );
  OAI21M1P U143 ( .A(n5), .B(n165), .C(n48), .Z(n256) );
  AOI22M1P U144 ( .A(n8), .B(\Queue[2][31] ), .C(\Queue[1][31] ), .D(n6), .Z(
        n51) );
  OAI21M1P U145 ( .A(n5), .B(n170), .C(n51), .Z(n281) );
  OAI21M1P U146 ( .A(n54), .B(n53), .C(n118), .Z(n55) );
  AOI21M1P U147 ( .A(n12), .B(n173), .C(n118), .Z(n80) );
  AOI22M1P U148 ( .A(\Queue[1][0] ), .B(n11), .C(n79), .D(Packet_Out[0]), .Z(
        n56) );
  OAI21M1P U149 ( .A(n121), .B(n82), .C(n56), .Z(n282) );
  AOI22M1P U150 ( .A(\Queue[1][1] ), .B(n11), .C(n79), .D(Packet_Out[1]), .Z(
        n57) );
  OAI21M1P U151 ( .A(n123), .B(n82), .C(n57), .Z(n283) );
  AOI22M1P U152 ( .A(\Queue[1][2] ), .B(n11), .C(n79), .D(Packet_Out[2]), .Z(
        n58) );
  OAI21M1P U153 ( .A(n125), .B(n82), .C(n58), .Z(n284) );
  AOI22M1P U154 ( .A(\Queue[1][3] ), .B(n11), .C(n79), .D(Packet_Out[3]), .Z(
        n59) );
  OAI21M1P U155 ( .A(n127), .B(n82), .C(n59), .Z(n285) );
  AOI22M1P U156 ( .A(\Queue[1][4] ), .B(n11), .C(n79), .D(Packet_Out[4]), .Z(
        n60) );
  OAI21M1P U157 ( .A(n129), .B(n82), .C(n60), .Z(n286) );
  AOI22M1P U158 ( .A(\Queue[1][5] ), .B(n11), .C(n79), .D(Packet_Out[5]), .Z(
        n61) );
  OAI21M1P U159 ( .A(n131), .B(n82), .C(n61), .Z(n287) );
  AOI22M1P U160 ( .A(\Queue[1][6] ), .B(n11), .C(n79), .D(Packet_Out[6]), .Z(
        n62) );
  OAI21M1P U161 ( .A(n133), .B(n82), .C(n62), .Z(n288) );
  AOI22M1P U162 ( .A(\Queue[1][7] ), .B(n11), .C(n79), .D(Packet_Out[7]), .Z(
        n63) );
  OAI21M1P U163 ( .A(n135), .B(n82), .C(n63), .Z(n298) );
  AOI22M1P U164 ( .A(\Queue[1][8] ), .B(n11), .C(n79), .D(Packet_Out[8]), .Z(
        n64) );
  OAI21M1P U165 ( .A(n137), .B(n82), .C(n64), .Z(n299) );
  AOI22M1P U166 ( .A(\Queue[1][9] ), .B(n11), .C(n79), .D(Packet_Out[9]), .Z(
        n65) );
  OAI21M1P U167 ( .A(n139), .B(n82), .C(n65), .Z(n300) );
  AOI22M1P U168 ( .A(\Queue[1][10] ), .B(n11), .C(n79), .D(Packet_Out[10]), 
        .Z(n66) );
  OAI21M1P U169 ( .A(n141), .B(n82), .C(n66), .Z(n301) );
  AOI22M1P U170 ( .A(\Queue[1][11] ), .B(n11), .C(n79), .D(Packet_Out[11]), 
        .Z(n67) );
  OAI21M1P U171 ( .A(n143), .B(n82), .C(n67), .Z(n302) );
  AOI22M1P U172 ( .A(\Queue[1][12] ), .B(n11), .C(n79), .D(Packet_Out[12]), 
        .Z(n68) );
  OAI21M1P U173 ( .A(n145), .B(n82), .C(n68), .Z(n303) );
  AOI22M1P U174 ( .A(\Queue[1][13] ), .B(n11), .C(n79), .D(Packet_Out[13]), 
        .Z(n69) );
  OAI21M1P U175 ( .A(n147), .B(n82), .C(n69), .Z(n304) );
  AOI22M1P U176 ( .A(\Queue[1][14] ), .B(n11), .C(n79), .D(Packet_Out[14]), 
        .Z(n70) );
  OAI21M1P U177 ( .A(n149), .B(n82), .C(n70), .Z(n305) );
  AOI22M1P U178 ( .A(\Queue[1][15] ), .B(n11), .C(n79), .D(Packet_Out[15]), 
        .Z(n71) );
  OAI21M1P U179 ( .A(n151), .B(n82), .C(n71), .Z(n306) );
  AOI22M1P U180 ( .A(\Queue[1][24] ), .B(n11), .C(n79), .D(Packet_Out[24]), 
        .Z(n72) );
  OAI21M1P U181 ( .A(n153), .B(n82), .C(n72), .Z(n307) );
  AOI22M1P U182 ( .A(\Queue[1][25] ), .B(n11), .C(n79), .D(Packet_Out[25]), 
        .Z(n73) );
  OAI21M1P U183 ( .A(n155), .B(n82), .C(n73), .Z(n308) );
  AOI22M1P U184 ( .A(\Queue[1][26] ), .B(n11), .C(n79), .D(Packet_Out[26]), 
        .Z(n74) );
  OAI21M1P U185 ( .A(n157), .B(n82), .C(n74), .Z(n309) );
  AOI22M1P U186 ( .A(\Queue[1][27] ), .B(n11), .C(n79), .D(Packet_Out[27]), 
        .Z(n75) );
  OAI21M1P U187 ( .A(n159), .B(n82), .C(n75), .Z(n310) );
  AOI22M1P U188 ( .A(\Queue[1][28] ), .B(n11), .C(n79), .D(Packet_Out[28]), 
        .Z(n76) );
  OAI21M1P U189 ( .A(n161), .B(n82), .C(n76), .Z(n311) );
  AOI22M1P U190 ( .A(\Queue[1][29] ), .B(n11), .C(n79), .D(Packet_Out[29]), 
        .Z(n77) );
  OAI21M1P U191 ( .A(n163), .B(n82), .C(n77), .Z(n312) );
  AOI22M1P U192 ( .A(\Queue[1][30] ), .B(n11), .C(n79), .D(Packet_Out[30]), 
        .Z(n78) );
  OAI21M1P U193 ( .A(n165), .B(n82), .C(n78), .Z(n313) );
  AOI22M1P U194 ( .A(\Queue[1][31] ), .B(n11), .C(n79), .D(Packet_Out[31]), 
        .Z(n81) );
  OAI21M1P U195 ( .A(n170), .B(n82), .C(n81), .Z(n314) );
  OA21M1P U196 ( .A(n116), .B(n85), .C(Rst_n), .Z(n83) );
  OAI211M1P U197 ( .A(n117), .B(n114), .C(n12), .D(n83), .Z(n112) );
  ND2M1P U198 ( .A(n84), .B(n114), .Z(n115) );
  AOI21M1P U199 ( .A(n12), .B(n117), .C(n118), .Z(n109) );
  AOI22M1P U200 ( .A(\Queue[2][0] ), .B(n7), .C(\Queue[3][0] ), .D(n9), .Z(n86) );
  OAI21M1P U201 ( .A(n121), .B(n3), .C(n86), .Z(n315) );
  AOI22M1P U202 ( .A(\Queue[2][1] ), .B(n7), .C(n9), .D(\Queue[3][1] ), .Z(n87) );
  OAI21M1P U203 ( .A(n123), .B(n3), .C(n87), .Z(n316) );
  AOI22M1P U204 ( .A(\Queue[2][2] ), .B(n7), .C(n9), .D(\Queue[3][2] ), .Z(n88) );
  OAI21M1P U205 ( .A(n125), .B(n3), .C(n88), .Z(n317) );
  AOI22M1P U206 ( .A(\Queue[2][3] ), .B(n7), .C(n9), .D(\Queue[3][3] ), .Z(n89) );
  OAI21M1P U207 ( .A(n127), .B(n3), .C(n89), .Z(n318) );
  AOI22M1P U208 ( .A(\Queue[2][4] ), .B(n7), .C(n9), .D(\Queue[3][4] ), .Z(n90) );
  OAI21M1P U209 ( .A(n129), .B(n3), .C(n90), .Z(n319) );
  AOI22M1P U210 ( .A(\Queue[2][5] ), .B(n7), .C(n9), .D(\Queue[3][5] ), .Z(n91) );
  OAI21M1P U211 ( .A(n131), .B(n3), .C(n91), .Z(n320) );
  AOI22M1P U212 ( .A(\Queue[2][6] ), .B(n7), .C(n9), .D(\Queue[3][6] ), .Z(n92) );
  OAI21M1P U213 ( .A(n133), .B(n3), .C(n92), .Z(n321) );
  AOI22M1P U214 ( .A(\Queue[2][7] ), .B(n7), .C(n9), .D(\Queue[3][7] ), .Z(n93) );
  OAI21M1P U215 ( .A(n135), .B(n3), .C(n93), .Z(n322) );
  AOI22M1P U216 ( .A(\Queue[2][8] ), .B(n7), .C(n9), .D(\Queue[3][8] ), .Z(n94) );
  OAI21M1P U217 ( .A(n137), .B(n3), .C(n94), .Z(n323) );
  AOI22M1P U218 ( .A(\Queue[2][9] ), .B(n7), .C(n9), .D(\Queue[3][9] ), .Z(n95) );
  OAI21M1P U219 ( .A(n139), .B(n3), .C(n95), .Z(n324) );
  AOI22M1P U220 ( .A(\Queue[2][10] ), .B(n7), .C(n9), .D(\Queue[3][10] ), .Z(
        n96) );
  OAI21M1P U221 ( .A(n141), .B(n3), .C(n96), .Z(n325) );
  AOI22M1P U222 ( .A(\Queue[2][11] ), .B(n7), .C(n9), .D(\Queue[3][11] ), .Z(
        n97) );
  OAI21M1P U223 ( .A(n143), .B(n3), .C(n97), .Z(n326) );
  AOI22M1P U224 ( .A(\Queue[2][12] ), .B(n7), .C(n9), .D(\Queue[3][12] ), .Z(
        n98) );
  OAI21M1P U225 ( .A(n145), .B(n3), .C(n98), .Z(n327) );
  AOI22M1P U226 ( .A(\Queue[2][13] ), .B(n7), .C(n9), .D(\Queue[3][13] ), .Z(
        n99) );
  OAI21M1P U227 ( .A(n147), .B(n3), .C(n99), .Z(n328) );
  AOI22M1P U228 ( .A(\Queue[2][14] ), .B(n7), .C(n9), .D(\Queue[3][14] ), .Z(
        n100) );
  OAI21M1P U229 ( .A(n149), .B(n3), .C(n100), .Z(n329) );
  AOI22M1P U230 ( .A(\Queue[2][15] ), .B(n7), .C(n9), .D(\Queue[3][15] ), .Z(
        n101) );
  OAI21M1P U231 ( .A(n151), .B(n3), .C(n101), .Z(n330) );
  AOI22M1P U232 ( .A(\Queue[2][24] ), .B(n7), .C(n9), .D(\Queue[3][24] ), .Z(
        n102) );
  OAI21M1P U233 ( .A(n153), .B(n3), .C(n102), .Z(n331) );
  AOI22M1P U234 ( .A(\Queue[2][25] ), .B(n7), .C(n9), .D(\Queue[3][25] ), .Z(
        n103) );
  OAI21M1P U235 ( .A(n155), .B(n3), .C(n103), .Z(n332) );
  AOI22M1P U236 ( .A(\Queue[2][26] ), .B(n7), .C(n9), .D(\Queue[3][26] ), .Z(
        n104) );
  OAI21M1P U237 ( .A(n157), .B(n3), .C(n104), .Z(n333) );
  AOI22M1P U238 ( .A(\Queue[2][27] ), .B(n7), .C(n9), .D(\Queue[3][27] ), .Z(
        n105) );
  OAI21M1P U239 ( .A(n159), .B(n3), .C(n105), .Z(n334) );
  AOI22M1P U240 ( .A(\Queue[2][28] ), .B(n7), .C(n9), .D(\Queue[3][28] ), .Z(
        n106) );
  OAI21M1P U241 ( .A(n161), .B(n3), .C(n106), .Z(n335) );
  AOI22M1P U242 ( .A(\Queue[2][29] ), .B(n7), .C(n9), .D(\Queue[3][29] ), .Z(
        n107) );
  OAI21M1P U243 ( .A(n163), .B(n3), .C(n107), .Z(n336) );
  AOI22M1P U244 ( .A(\Queue[2][30] ), .B(n7), .C(n9), .D(\Queue[3][30] ), .Z(
        n108) );
  OAI21M1P U245 ( .A(n165), .B(n3), .C(n108), .Z(n337) );
  AOI22M1P U246 ( .A(\Queue[2][31] ), .B(n7), .C(n9), .D(\Queue[3][31] ), .Z(
        n111) );
  OAI21M1P U247 ( .A(n170), .B(n3), .C(n111), .Z(n338) );
  OA21M1P U248 ( .A(n116), .B(n117), .C(Rst_n), .Z(n113) );
  OAI211M1P U249 ( .A(n119), .B(n114), .C(n12), .D(n113), .Z(n169) );
  AOI21M1P U250 ( .A(n12), .B(n119), .C(n118), .Z(n166) );
  AOI22M1P U251 ( .A(\Queue[3][0] ), .B(n13), .C(n10), .D(\Queue[4][0] ), .Z(
        n120) );
  OAI21M1P U252 ( .A(n121), .B(n4), .C(n120), .Z(n339) );
  AOI22M1P U253 ( .A(\Queue[3][1] ), .B(n13), .C(n10), .D(\Queue[4][1] ), .Z(
        n122) );
  OAI21M1P U254 ( .A(n123), .B(n4), .C(n122), .Z(n340) );
  AOI22M1P U255 ( .A(\Queue[3][2] ), .B(n13), .C(n10), .D(\Queue[4][2] ), .Z(
        n124) );
  OAI21M1P U256 ( .A(n125), .B(n4), .C(n124), .Z(n341) );
  AOI22M1P U257 ( .A(\Queue[3][3] ), .B(n13), .C(n10), .D(\Queue[4][3] ), .Z(
        n126) );
  OAI21M1P U258 ( .A(n127), .B(n4), .C(n126), .Z(n342) );
  AOI22M1P U259 ( .A(\Queue[3][4] ), .B(n13), .C(n10), .D(\Queue[4][4] ), .Z(
        n128) );
  OAI21M1P U260 ( .A(n129), .B(n4), .C(n128), .Z(n343) );
  AOI22M1P U261 ( .A(\Queue[3][5] ), .B(n13), .C(n10), .D(\Queue[4][5] ), .Z(
        n130) );
  OAI21M1P U262 ( .A(n131), .B(n4), .C(n130), .Z(n344) );
  AOI22M1P U263 ( .A(\Queue[3][6] ), .B(n13), .C(n10), .D(\Queue[4][6] ), .Z(
        n132) );
  OAI21M1P U264 ( .A(n133), .B(n4), .C(n132), .Z(n345) );
  AOI22M1P U265 ( .A(\Queue[3][7] ), .B(n13), .C(n10), .D(\Queue[4][7] ), .Z(
        n134) );
  OAI21M1P U266 ( .A(n135), .B(n4), .C(n134), .Z(n346) );
  AOI22M1P U267 ( .A(\Queue[3][8] ), .B(n13), .C(n10), .D(\Queue[4][8] ), .Z(
        n136) );
  OAI21M1P U268 ( .A(n137), .B(n4), .C(n136), .Z(n347) );
  AOI22M1P U269 ( .A(\Queue[3][9] ), .B(n13), .C(n10), .D(\Queue[4][9] ), .Z(
        n138) );
  OAI21M1P U270 ( .A(n139), .B(n4), .C(n138), .Z(n348) );
  AOI22M1P U271 ( .A(\Queue[3][10] ), .B(n13), .C(n10), .D(\Queue[4][10] ), 
        .Z(n140) );
  OAI21M1P U272 ( .A(n141), .B(n4), .C(n140), .Z(n349) );
  AOI22M1P U273 ( .A(\Queue[3][11] ), .B(n13), .C(n10), .D(\Queue[4][11] ), 
        .Z(n142) );
  OAI21M1P U274 ( .A(n143), .B(n4), .C(n142), .Z(n350) );
  AOI22M1P U275 ( .A(\Queue[3][12] ), .B(n13), .C(n10), .D(\Queue[4][12] ), 
        .Z(n144) );
  OAI21M1P U276 ( .A(n145), .B(n4), .C(n144), .Z(n351) );
  AOI22M1P U277 ( .A(\Queue[3][13] ), .B(n13), .C(n10), .D(\Queue[4][13] ), 
        .Z(n146) );
  OAI21M1P U278 ( .A(n147), .B(n4), .C(n146), .Z(n352) );
  AOI22M1P U279 ( .A(\Queue[3][14] ), .B(n13), .C(n10), .D(\Queue[4][14] ), 
        .Z(n148) );
  OAI21M1P U280 ( .A(n149), .B(n4), .C(n148), .Z(n353) );
  AOI22M1P U281 ( .A(\Queue[3][15] ), .B(n13), .C(n10), .D(\Queue[4][15] ), 
        .Z(n150) );
  OAI21M1P U282 ( .A(n151), .B(n4), .C(n150), .Z(n354) );
  AOI22M1P U283 ( .A(\Queue[3][24] ), .B(n13), .C(n10), .D(\Queue[4][24] ), 
        .Z(n152) );
  OAI21M1P U284 ( .A(n153), .B(n4), .C(n152), .Z(n355) );
  AOI22M1P U285 ( .A(\Queue[3][25] ), .B(n13), .C(n10), .D(\Queue[4][25] ), 
        .Z(n154) );
  OAI21M1P U286 ( .A(n155), .B(n4), .C(n154), .Z(n356) );
  AOI22M1P U287 ( .A(\Queue[3][26] ), .B(n13), .C(n10), .D(\Queue[4][26] ), 
        .Z(n156) );
  OAI21M1P U288 ( .A(n157), .B(n4), .C(n156), .Z(n357) );
  AOI22M1P U289 ( .A(\Queue[3][27] ), .B(n13), .C(n10), .D(\Queue[4][27] ), 
        .Z(n158) );
  OAI21M1P U290 ( .A(n159), .B(n4), .C(n158), .Z(n358) );
  AOI22M1P U291 ( .A(\Queue[3][28] ), .B(n167), .C(n10), .D(\Queue[4][28] ), 
        .Z(n160) );
  OAI21M1P U292 ( .A(n161), .B(n4), .C(n160), .Z(n359) );
  AOI22M1P U293 ( .A(\Queue[3][29] ), .B(n167), .C(n10), .D(\Queue[4][29] ), 
        .Z(n162) );
  OAI21M1P U294 ( .A(n163), .B(n4), .C(n162), .Z(n360) );
  AOI22M1P U295 ( .A(\Queue[3][30] ), .B(n167), .C(n10), .D(\Queue[4][30] ), 
        .Z(n164) );
  OAI21M1P U296 ( .A(n165), .B(n4), .C(n164), .Z(n361) );
  AOI22M1P U297 ( .A(\Queue[3][31] ), .B(n13), .C(n10), .D(\Queue[4][31] ), 
        .Z(n168) );
  OAI21M1P U298 ( .A(n170), .B(n4), .C(n168), .Z(n362) );
  AOI22M1P U299 ( .A(n173), .B(n172), .C(n171), .D(Empty), .Z(n364) );
endmodule


module Node_Manager ( Clk_r, Rst_n, Packet_From_Core, Packet_From_Node, 
        Packet_From_Node_Valid, Read_Packet, To_Node_Write, Router_Address, 
        Link_Config, Packet_To_Core, Packet_To_Node, Packet_To_Node_Valid, 
        Core_Load_Ack, Queue_Empty, To_Node_Full );
  input [31:0] Packet_From_Core;
  input [31:0] Packet_From_Node;
  output [7:0] Router_Address;
  output [3:0] Link_Config;
  output [31:0] Packet_To_Core;
  output [31:0] Packet_To_Node;
  input Clk_r, Rst_n, Packet_From_Node_Valid, Read_Packet, To_Node_Write;
  output Packet_To_Node_Valid, Core_Load_Ack, Queue_Empty, To_Node_Full;
  wire   Write_Queue, Queue_Full, Read_Out_Queue, Out_Queue_Empty, N8, N42,
         N43, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7;

  Packet_Queue_2 In_Queue ( .Clk_r(Clk_r), .Rst_n(Rst_n), .Packet_In({
        Packet_From_Node[31:24], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, Packet_From_Node[15:0]}), .Read_Ack(Read_Packet), .Write_Ack(
        Write_Queue), .Packet_Out({Packet_To_Core[31:24], 
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, Packet_To_Core[15:0]}), .Empty(Queue_Empty), .Full(Queue_Full) );
  Packet_Queue_1 Out_Queue ( .Clk_r(Clk_r), .Rst_n(Rst_n), .Packet_In(
        Packet_From_Core), .Read_Ack(Read_Out_Queue), .Write_Ack(To_Node_Write), .Packet_Out(Packet_To_Node), .Empty(Out_Queue_Empty), .Full(To_Node_Full) );
  FD2LQM1P \Router_Address_reg[0]  ( .D(Packet_From_Node[0]), .LD(n2), .CP(
        Clk_r), .CD(Rst_n), .Q(Router_Address[0]) );
  FD2LQM1P \Router_Address_reg[1]  ( .D(Packet_From_Node[1]), .LD(n2), .CP(
        Clk_r), .CD(Rst_n), .Q(Router_Address[1]) );
  FD2LQM1P \Router_Address_reg[2]  ( .D(Packet_From_Node[2]), .LD(n2), .CP(
        Clk_r), .CD(Rst_n), .Q(Router_Address[2]) );
  FD2LQM1P \Router_Address_reg[3]  ( .D(Packet_From_Node[3]), .LD(n2), .CP(
        Clk_r), .CD(Rst_n), .Q(Router_Address[3]) );
  FD2LQM1P \Router_Address_reg[4]  ( .D(Packet_From_Node[4]), .LD(n2), .CP(
        Clk_r), .CD(Rst_n), .Q(Router_Address[4]) );
  FD2LQM1P \Router_Address_reg[5]  ( .D(Packet_From_Node[5]), .LD(n2), .CP(
        Clk_r), .CD(Rst_n), .Q(Router_Address[5]) );
  FD2LQM1P \Router_Address_reg[6]  ( .D(Packet_From_Node[6]), .LD(n2), .CP(
        Clk_r), .CD(Rst_n), .Q(Router_Address[6]) );
  FD2LQM1P \Router_Address_reg[7]  ( .D(Packet_From_Node[7]), .LD(n2), .CP(
        Clk_r), .CD(Rst_n), .Q(Router_Address[7]) );
  FD2LQM1P \Link_Config_reg[0]  ( .D(Packet_From_Node[0]), .LD(n1), .CP(Clk_r), 
        .CD(Rst_n), .Q(Link_Config[0]) );
  FD2LQM1P \Link_Config_reg[1]  ( .D(Packet_From_Node[1]), .LD(n1), .CP(Clk_r), 
        .CD(Rst_n), .Q(Link_Config[1]) );
  FD2LQM1P \Link_Config_reg[2]  ( .D(Packet_From_Node[2]), .LD(n1), .CP(Clk_r), 
        .CD(Rst_n), .Q(Link_Config[2]) );
  FD2LQM1P \Link_Config_reg[3]  ( .D(Packet_From_Node[3]), .LD(n1), .CP(Clk_r), 
        .CD(Rst_n), .Q(Link_Config[3]) );
  FD2QM1P Read_Out_Queue_reg ( .D(Packet_To_Node_Valid), .CP(Clk_r), .CD(Rst_n), .Q(Read_Out_Queue) );
  FD2QM1P Packet_To_Node_Valid_reg ( .D(N8), .CP(Clk_r), .CD(Rst_n), .Q(
        Packet_To_Node_Valid) );
  FD2QM1P Core_Load_Ack_reg ( .D(N42), .CP(Clk_r), .CD(Rst_n), .Q(
        Core_Load_Ack) );
  FD2QM1P Write_Queue_reg ( .D(N43), .CP(Clk_r), .CD(Rst_n), .Q(Write_Queue)
         );
  NR2M1P U3 ( .A(Packet_From_Node[16]), .B(n10), .Z(n2) );
  ND4M1P U5 ( .A(Packet_From_Node[30]), .B(Packet_From_Node[31]), .C(
        Packet_From_Node[28]), .D(Packet_From_Node[29]), .Z(n5) );
  ND4M1P U6 ( .A(Packet_From_Node[26]), .B(Packet_From_Node[27]), .C(
        Packet_From_Node[24]), .D(Packet_From_Node[25]), .Z(n4) );
  AND2M1P U7 ( .A(n5), .B(n4), .Z(n3) );
  ND2BNM1P U8 ( .B(Core_Load_Ack), .A(Packet_From_Node_Valid), .Z(n6) );
  AOI21M1P U9 ( .A(n3), .B(Queue_Full), .C(n6), .Z(N42) );
  NR3CNM1P U10 ( .C(n3), .A(Queue_Full), .B(n6), .Z(N43) );
  NR2M1P U11 ( .A(Out_Queue_Empty), .B(Packet_To_Node_Valid), .Z(N8) );
  NR3M1P U12 ( .A(Packet_From_Node[23]), .B(Packet_From_Node[18]), .C(
        Packet_From_Node[17]), .Z(n9) );
  NR3M1P U13 ( .A(Packet_From_Node[19]), .B(Packet_From_Node[20]), .C(n4), .Z(
        n8) );
  NR3M1P U14 ( .A(Packet_From_Node[21]), .B(n6), .C(n5), .Z(n7) );
  ND4DNM1P U15 ( .D(Packet_From_Node[22]), .A(n9), .B(n8), .C(n7), .Z(n10) );
  NR2BNM1P U16 ( .B(Packet_From_Node[16]), .A(n10), .Z(n1) );
endmodule


module Packet_Queue_3 ( Clk_r, Rst_n, Packet_In, Read_Ack, Write_Ack, 
        Packet_Out, Empty, Full );
  input [31:0] Packet_In;
  output [31:0] Packet_Out;
  input Clk_r, Rst_n, Read_Ack, Write_Ack;
  output Empty, Full;
  wire   \Queue[4][31] , \Queue[4][30] , \Queue[4][29] , \Queue[4][28] ,
         \Queue[4][27] , \Queue[4][26] , \Queue[4][25] , \Queue[4][24] ,
         \Queue[4][23] , \Queue[4][22] , \Queue[4][21] , \Queue[4][20] ,
         \Queue[4][19] , \Queue[4][18] , \Queue[4][17] , \Queue[4][16] ,
         \Queue[4][15] , \Queue[4][14] , \Queue[4][13] , \Queue[4][12] ,
         \Queue[4][11] , \Queue[4][10] , \Queue[4][9] , \Queue[4][8] ,
         \Queue[4][7] , \Queue[4][6] , \Queue[4][5] , \Queue[4][4] ,
         \Queue[4][3] , \Queue[4][2] , \Queue[4][1] , \Queue[4][0] ,
         \Queue[3][31] , \Queue[3][30] , \Queue[3][29] , \Queue[3][28] ,
         \Queue[3][27] , \Queue[3][26] , \Queue[3][25] , \Queue[3][24] ,
         \Queue[3][23] , \Queue[3][22] , \Queue[3][21] , \Queue[3][20] ,
         \Queue[3][19] , \Queue[3][18] , \Queue[3][17] , \Queue[3][16] ,
         \Queue[3][15] , \Queue[3][14] , \Queue[3][13] , \Queue[3][12] ,
         \Queue[3][11] , \Queue[3][10] , \Queue[3][9] , \Queue[3][8] ,
         \Queue[3][7] , \Queue[3][6] , \Queue[3][5] , \Queue[3][4] ,
         \Queue[3][3] , \Queue[3][2] , \Queue[3][1] , \Queue[3][0] ,
         \Queue[2][31] , \Queue[2][30] , \Queue[2][29] , \Queue[2][28] ,
         \Queue[2][27] , \Queue[2][26] , \Queue[2][25] , \Queue[2][24] ,
         \Queue[2][23] , \Queue[2][22] , \Queue[2][21] , \Queue[2][20] ,
         \Queue[2][19] , \Queue[2][18] , \Queue[2][17] , \Queue[2][16] ,
         \Queue[2][15] , \Queue[2][14] , \Queue[2][13] , \Queue[2][12] ,
         \Queue[2][11] , \Queue[2][10] , \Queue[2][9] , \Queue[2][8] ,
         \Queue[2][7] , \Queue[2][6] , \Queue[2][5] , \Queue[2][4] ,
         \Queue[2][3] , \Queue[2][2] , \Queue[2][1] , \Queue[2][0] ,
         \Queue[1][31] , \Queue[1][30] , \Queue[1][29] , \Queue[1][28] ,
         \Queue[1][27] , \Queue[1][26] , \Queue[1][25] , \Queue[1][24] ,
         \Queue[1][23] , \Queue[1][22] , \Queue[1][21] , \Queue[1][20] ,
         \Queue[1][19] , \Queue[1][18] , \Queue[1][17] , \Queue[1][16] ,
         \Queue[1][15] , \Queue[1][14] , \Queue[1][13] , \Queue[1][12] ,
         \Queue[1][11] , \Queue[1][10] , \Queue[1][9] , \Queue[1][8] ,
         \Queue[1][7] , \Queue[1][6] , \Queue[1][5] , \Queue[1][4] ,
         \Queue[1][3] , \Queue[1][2] , \Queue[1][1] , \Queue[1][0] , n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542;
  wire   [2:0] Count;

  FDN2QM1P \Count_reg[0]  ( .D(n377), .CPN(Clk_r), .CD(Rst_n), .Q(Count[0]) );
  FDN2QM1P \Count_reg[1]  ( .D(n378), .CPN(Clk_r), .CD(Rst_n), .Q(Count[1]) );
  FDN2QM1P \Count_reg[2]  ( .D(n379), .CPN(Clk_r), .CD(Rst_n), .Q(Count[2]) );
  FDN1QM1P \Queue_reg[4][30]  ( .D(n411), .CPN(Clk_r), .Q(\Queue[4][30] ) );
  FDN1QM1P \Queue_reg[3][30]  ( .D(n539), .CPN(Clk_r), .Q(\Queue[3][30] ) );
  FDN1QM1P \Queue_reg[2][30]  ( .D(n507), .CPN(Clk_r), .Q(\Queue[2][30] ) );
  FDN1QM1P \Queue_reg[4][29]  ( .D(n410), .CPN(Clk_r), .Q(\Queue[4][29] ) );
  FDN1QM1P \Queue_reg[3][29]  ( .D(n538), .CPN(Clk_r), .Q(\Queue[3][29] ) );
  FDN1QM1P \Queue_reg[2][29]  ( .D(n506), .CPN(Clk_r), .Q(\Queue[2][29] ) );
  FDN1QM1P \Queue_reg[4][28]  ( .D(n409), .CPN(Clk_r), .Q(\Queue[4][28] ) );
  FDN1QM1P \Queue_reg[3][28]  ( .D(n537), .CPN(Clk_r), .Q(\Queue[3][28] ) );
  FDN1QM1P \Queue_reg[2][28]  ( .D(n505), .CPN(Clk_r), .Q(\Queue[2][28] ) );
  FDN1QM1P \Queue_reg[4][27]  ( .D(n408), .CPN(Clk_r), .Q(\Queue[4][27] ) );
  FDN1QM1P \Queue_reg[3][27]  ( .D(n536), .CPN(Clk_r), .Q(\Queue[3][27] ) );
  FDN1QM1P \Queue_reg[2][27]  ( .D(n504), .CPN(Clk_r), .Q(\Queue[2][27] ) );
  FDN1QM1P \Queue_reg[4][26]  ( .D(n407), .CPN(Clk_r), .Q(\Queue[4][26] ) );
  FDN1QM1P \Queue_reg[3][26]  ( .D(n535), .CPN(Clk_r), .Q(\Queue[3][26] ) );
  FDN1QM1P \Queue_reg[2][26]  ( .D(n503), .CPN(Clk_r), .Q(\Queue[2][26] ) );
  FDN1QM1P \Queue_reg[4][25]  ( .D(n406), .CPN(Clk_r), .Q(\Queue[4][25] ) );
  FDN1QM1P \Queue_reg[3][25]  ( .D(n534), .CPN(Clk_r), .Q(\Queue[3][25] ) );
  FDN1QM1P \Queue_reg[2][25]  ( .D(n502), .CPN(Clk_r), .Q(\Queue[2][25] ) );
  FDN1QM1P \Queue_reg[4][24]  ( .D(n405), .CPN(Clk_r), .Q(\Queue[4][24] ) );
  FDN1QM1P \Queue_reg[3][24]  ( .D(n533), .CPN(Clk_r), .Q(\Queue[3][24] ) );
  FDN1QM1P \Queue_reg[2][24]  ( .D(n501), .CPN(Clk_r), .Q(\Queue[2][24] ) );
  FDN1QM1P \Queue_reg[4][23]  ( .D(n404), .CPN(Clk_r), .Q(\Queue[4][23] ) );
  FDN1QM1P \Queue_reg[3][23]  ( .D(n532), .CPN(Clk_r), .Q(\Queue[3][23] ) );
  FDN1QM1P \Queue_reg[2][23]  ( .D(n500), .CPN(Clk_r), .Q(\Queue[2][23] ) );
  FDN1QM1P \Queue_reg[4][22]  ( .D(n403), .CPN(Clk_r), .Q(\Queue[4][22] ) );
  FDN1QM1P \Queue_reg[3][22]  ( .D(n531), .CPN(Clk_r), .Q(\Queue[3][22] ) );
  FDN1QM1P \Queue_reg[2][22]  ( .D(n499), .CPN(Clk_r), .Q(\Queue[2][22] ) );
  FDN1QM1P \Queue_reg[4][21]  ( .D(n402), .CPN(Clk_r), .Q(\Queue[4][21] ) );
  FDN1QM1P \Queue_reg[3][21]  ( .D(n530), .CPN(Clk_r), .Q(\Queue[3][21] ) );
  FDN1QM1P \Queue_reg[2][21]  ( .D(n498), .CPN(Clk_r), .Q(\Queue[2][21] ) );
  FDN1QM1P \Queue_reg[4][20]  ( .D(n401), .CPN(Clk_r), .Q(\Queue[4][20] ) );
  FDN1QM1P \Queue_reg[3][20]  ( .D(n529), .CPN(Clk_r), .Q(\Queue[3][20] ) );
  FDN1QM1P \Queue_reg[2][20]  ( .D(n497), .CPN(Clk_r), .Q(\Queue[2][20] ) );
  FDN1QM1P \Queue_reg[4][19]  ( .D(n400), .CPN(Clk_r), .Q(\Queue[4][19] ) );
  FDN1QM1P \Queue_reg[3][19]  ( .D(n528), .CPN(Clk_r), .Q(\Queue[3][19] ) );
  FDN1QM1P \Queue_reg[2][19]  ( .D(n496), .CPN(Clk_r), .Q(\Queue[2][19] ) );
  FDN1QM1P \Queue_reg[4][18]  ( .D(n399), .CPN(Clk_r), .Q(\Queue[4][18] ) );
  FDN1QM1P \Queue_reg[3][18]  ( .D(n527), .CPN(Clk_r), .Q(\Queue[3][18] ) );
  FDN1QM1P \Queue_reg[2][18]  ( .D(n495), .CPN(Clk_r), .Q(\Queue[2][18] ) );
  FDN1QM1P \Queue_reg[4][17]  ( .D(n398), .CPN(Clk_r), .Q(\Queue[4][17] ) );
  FDN1QM1P \Queue_reg[3][17]  ( .D(n526), .CPN(Clk_r), .Q(\Queue[3][17] ) );
  FDN1QM1P \Queue_reg[2][17]  ( .D(n494), .CPN(Clk_r), .Q(\Queue[2][17] ) );
  FDN1QM1P \Queue_reg[4][16]  ( .D(n397), .CPN(Clk_r), .Q(\Queue[4][16] ) );
  FDN1QM1P \Queue_reg[3][16]  ( .D(n525), .CPN(Clk_r), .Q(\Queue[3][16] ) );
  FDN1QM1P \Queue_reg[2][16]  ( .D(n493), .CPN(Clk_r), .Q(\Queue[2][16] ) );
  FDN1QM1P \Queue_reg[4][15]  ( .D(n396), .CPN(Clk_r), .Q(\Queue[4][15] ) );
  FDN1QM1P \Queue_reg[3][15]  ( .D(n524), .CPN(Clk_r), .Q(\Queue[3][15] ) );
  FDN1QM1P \Queue_reg[2][15]  ( .D(n492), .CPN(Clk_r), .Q(\Queue[2][15] ) );
  FDN1QM1P \Queue_reg[4][14]  ( .D(n395), .CPN(Clk_r), .Q(\Queue[4][14] ) );
  FDN1QM1P \Queue_reg[3][14]  ( .D(n523), .CPN(Clk_r), .Q(\Queue[3][14] ) );
  FDN1QM1P \Queue_reg[2][14]  ( .D(n491), .CPN(Clk_r), .Q(\Queue[2][14] ) );
  FDN1QM1P \Queue_reg[4][13]  ( .D(n394), .CPN(Clk_r), .Q(\Queue[4][13] ) );
  FDN1QM1P \Queue_reg[3][13]  ( .D(n522), .CPN(Clk_r), .Q(\Queue[3][13] ) );
  FDN1QM1P \Queue_reg[2][13]  ( .D(n490), .CPN(Clk_r), .Q(\Queue[2][13] ) );
  FDN1QM1P \Queue_reg[4][12]  ( .D(n393), .CPN(Clk_r), .Q(\Queue[4][12] ) );
  FDN1QM1P \Queue_reg[3][12]  ( .D(n521), .CPN(Clk_r), .Q(\Queue[3][12] ) );
  FDN1QM1P \Queue_reg[2][12]  ( .D(n489), .CPN(Clk_r), .Q(\Queue[2][12] ) );
  FDN1QM1P \Queue_reg[4][11]  ( .D(n392), .CPN(Clk_r), .Q(\Queue[4][11] ) );
  FDN1QM1P \Queue_reg[3][11]  ( .D(n520), .CPN(Clk_r), .Q(\Queue[3][11] ) );
  FDN1QM1P \Queue_reg[2][11]  ( .D(n488), .CPN(Clk_r), .Q(\Queue[2][11] ) );
  FDN1QM1P \Queue_reg[4][10]  ( .D(n391), .CPN(Clk_r), .Q(\Queue[4][10] ) );
  FDN1QM1P \Queue_reg[3][10]  ( .D(n519), .CPN(Clk_r), .Q(\Queue[3][10] ) );
  FDN1QM1P \Queue_reg[2][10]  ( .D(n487), .CPN(Clk_r), .Q(\Queue[2][10] ) );
  FDN1QM1P \Queue_reg[4][9]  ( .D(n390), .CPN(Clk_r), .Q(\Queue[4][9] ) );
  FDN1QM1P \Queue_reg[3][9]  ( .D(n518), .CPN(Clk_r), .Q(\Queue[3][9] ) );
  FDN1QM1P \Queue_reg[2][9]  ( .D(n486), .CPN(Clk_r), .Q(\Queue[2][9] ) );
  FDN1QM1P \Queue_reg[4][8]  ( .D(n389), .CPN(Clk_r), .Q(\Queue[4][8] ) );
  FDN1QM1P \Queue_reg[3][8]  ( .D(n517), .CPN(Clk_r), .Q(\Queue[3][8] ) );
  FDN1QM1P \Queue_reg[2][8]  ( .D(n485), .CPN(Clk_r), .Q(\Queue[2][8] ) );
  FDN1QM1P \Queue_reg[4][7]  ( .D(n388), .CPN(Clk_r), .Q(\Queue[4][7] ) );
  FDN1QM1P \Queue_reg[3][7]  ( .D(n516), .CPN(Clk_r), .Q(\Queue[3][7] ) );
  FDN1QM1P \Queue_reg[2][7]  ( .D(n484), .CPN(Clk_r), .Q(\Queue[2][7] ) );
  FDN1QM1P \Queue_reg[4][6]  ( .D(n387), .CPN(Clk_r), .Q(\Queue[4][6] ) );
  FDN1QM1P \Queue_reg[3][6]  ( .D(n515), .CPN(Clk_r), .Q(\Queue[3][6] ) );
  FDN1QM1P \Queue_reg[2][6]  ( .D(n483), .CPN(Clk_r), .Q(\Queue[2][6] ) );
  FDN1QM1P \Queue_reg[4][5]  ( .D(n386), .CPN(Clk_r), .Q(\Queue[4][5] ) );
  FDN1QM1P \Queue_reg[3][5]  ( .D(n514), .CPN(Clk_r), .Q(\Queue[3][5] ) );
  FDN1QM1P \Queue_reg[2][5]  ( .D(n482), .CPN(Clk_r), .Q(\Queue[2][5] ) );
  FDN1QM1P \Queue_reg[4][4]  ( .D(n385), .CPN(Clk_r), .Q(\Queue[4][4] ) );
  FDN1QM1P \Queue_reg[3][4]  ( .D(n513), .CPN(Clk_r), .Q(\Queue[3][4] ) );
  FDN1QM1P \Queue_reg[2][4]  ( .D(n481), .CPN(Clk_r), .Q(\Queue[2][4] ) );
  FDN1QM1P \Queue_reg[4][3]  ( .D(n384), .CPN(Clk_r), .Q(\Queue[4][3] ) );
  FDN1QM1P \Queue_reg[3][3]  ( .D(n512), .CPN(Clk_r), .Q(\Queue[3][3] ) );
  FDN1QM1P \Queue_reg[2][3]  ( .D(n480), .CPN(Clk_r), .Q(\Queue[2][3] ) );
  FDN1QM1P \Queue_reg[4][2]  ( .D(n383), .CPN(Clk_r), .Q(\Queue[4][2] ) );
  FDN1QM1P \Queue_reg[3][2]  ( .D(n511), .CPN(Clk_r), .Q(\Queue[3][2] ) );
  FDN1QM1P \Queue_reg[2][2]  ( .D(n479), .CPN(Clk_r), .Q(\Queue[2][2] ) );
  FDN1QM1P \Queue_reg[4][1]  ( .D(n382), .CPN(Clk_r), .Q(\Queue[4][1] ) );
  FDN1QM1P \Queue_reg[3][1]  ( .D(n510), .CPN(Clk_r), .Q(\Queue[3][1] ) );
  FDN1QM1P \Queue_reg[2][1]  ( .D(n478), .CPN(Clk_r), .Q(\Queue[2][1] ) );
  FDN1QM1P \Queue_reg[4][0]  ( .D(n381), .CPN(Clk_r), .Q(\Queue[4][0] ) );
  FDN1QM1P \Queue_reg[3][0]  ( .D(n509), .CPN(Clk_r), .Q(\Queue[3][0] ) );
  FDN1QM1P \Queue_reg[2][0]  ( .D(n477), .CPN(Clk_r), .Q(\Queue[2][0] ) );
  FDN1QM1P \Queue_reg[4][31]  ( .D(n380), .CPN(Clk_r), .Q(\Queue[4][31] ) );
  FDN1QM1P \Queue_reg[3][31]  ( .D(n540), .CPN(Clk_r), .Q(\Queue[3][31] ) );
  FDN1QM1P \Queue_reg[2][31]  ( .D(n508), .CPN(Clk_r), .Q(\Queue[2][31] ) );
  FDN2QM1P Full_reg ( .D(n412), .CPN(Clk_r), .CD(Rst_n), .Q(Full) );
  FDN1QM1P \Queue_reg[1][31]  ( .D(n444), .CPN(Clk_r), .Q(\Queue[1][31] ) );
  FDN1QM1P \Queue_reg[0][31]  ( .D(n476), .CPN(Clk_r), .Q(Packet_Out[31]) );
  FDN1QM1P \Queue_reg[1][30]  ( .D(n443), .CPN(Clk_r), .Q(\Queue[1][30] ) );
  FDN1QM1P \Queue_reg[0][30]  ( .D(n475), .CPN(Clk_r), .Q(Packet_Out[30]) );
  FDN1QM1P \Queue_reg[1][29]  ( .D(n442), .CPN(Clk_r), .Q(\Queue[1][29] ) );
  FDN1QM1P \Queue_reg[0][29]  ( .D(n474), .CPN(Clk_r), .Q(Packet_Out[29]) );
  FDN1QM1P \Queue_reg[1][28]  ( .D(n441), .CPN(Clk_r), .Q(\Queue[1][28] ) );
  FDN1QM1P \Queue_reg[0][28]  ( .D(n473), .CPN(Clk_r), .Q(Packet_Out[28]) );
  FDN1QM1P \Queue_reg[1][27]  ( .D(n440), .CPN(Clk_r), .Q(\Queue[1][27] ) );
  FDN1QM1P \Queue_reg[0][27]  ( .D(n472), .CPN(Clk_r), .Q(Packet_Out[27]) );
  FDN1QM1P \Queue_reg[1][26]  ( .D(n439), .CPN(Clk_r), .Q(\Queue[1][26] ) );
  FDN1QM1P \Queue_reg[0][26]  ( .D(n471), .CPN(Clk_r), .Q(Packet_Out[26]) );
  FDN1QM1P \Queue_reg[1][25]  ( .D(n438), .CPN(Clk_r), .Q(\Queue[1][25] ) );
  FDN1QM1P \Queue_reg[0][25]  ( .D(n470), .CPN(Clk_r), .Q(Packet_Out[25]) );
  FDN1QM1P \Queue_reg[1][24]  ( .D(n437), .CPN(Clk_r), .Q(\Queue[1][24] ) );
  FDN1QM1P \Queue_reg[0][24]  ( .D(n469), .CPN(Clk_r), .Q(Packet_Out[24]) );
  FDN1QM1P \Queue_reg[1][23]  ( .D(n436), .CPN(Clk_r), .Q(\Queue[1][23] ) );
  FDN1QM1P \Queue_reg[0][23]  ( .D(n468), .CPN(Clk_r), .Q(Packet_Out[23]) );
  FDN1QM1P \Queue_reg[1][22]  ( .D(n435), .CPN(Clk_r), .Q(\Queue[1][22] ) );
  FDN1QM1P \Queue_reg[0][22]  ( .D(n467), .CPN(Clk_r), .Q(Packet_Out[22]) );
  FDN1QM1P \Queue_reg[1][21]  ( .D(n434), .CPN(Clk_r), .Q(\Queue[1][21] ) );
  FDN1QM1P \Queue_reg[0][21]  ( .D(n466), .CPN(Clk_r), .Q(Packet_Out[21]) );
  FDN1QM1P \Queue_reg[1][20]  ( .D(n433), .CPN(Clk_r), .Q(\Queue[1][20] ) );
  FDN1QM1P \Queue_reg[0][20]  ( .D(n465), .CPN(Clk_r), .Q(Packet_Out[20]) );
  FDN1QM1P \Queue_reg[1][19]  ( .D(n432), .CPN(Clk_r), .Q(\Queue[1][19] ) );
  FDN1QM1P \Queue_reg[0][19]  ( .D(n464), .CPN(Clk_r), .Q(Packet_Out[19]) );
  FDN1QM1P \Queue_reg[1][18]  ( .D(n431), .CPN(Clk_r), .Q(\Queue[1][18] ) );
  FDN1QM1P \Queue_reg[0][18]  ( .D(n463), .CPN(Clk_r), .Q(Packet_Out[18]) );
  FDN1QM1P \Queue_reg[1][17]  ( .D(n430), .CPN(Clk_r), .Q(\Queue[1][17] ) );
  FDN1QM1P \Queue_reg[0][17]  ( .D(n462), .CPN(Clk_r), .Q(Packet_Out[17]) );
  FDN1QM1P \Queue_reg[1][16]  ( .D(n429), .CPN(Clk_r), .Q(\Queue[1][16] ) );
  FDN1QM1P \Queue_reg[0][16]  ( .D(n461), .CPN(Clk_r), .Q(Packet_Out[16]) );
  FDN1QM1P \Queue_reg[1][15]  ( .D(n428), .CPN(Clk_r), .Q(\Queue[1][15] ) );
  FDN1QM1P \Queue_reg[0][15]  ( .D(n460), .CPN(Clk_r), .Q(Packet_Out[15]) );
  FDN1QM1P \Queue_reg[1][14]  ( .D(n427), .CPN(Clk_r), .Q(\Queue[1][14] ) );
  FDN1QM1P \Queue_reg[0][14]  ( .D(n459), .CPN(Clk_r), .Q(Packet_Out[14]) );
  FDN1QM1P \Queue_reg[1][13]  ( .D(n426), .CPN(Clk_r), .Q(\Queue[1][13] ) );
  FDN1QM1P \Queue_reg[0][13]  ( .D(n458), .CPN(Clk_r), .Q(Packet_Out[13]) );
  FDN1QM1P \Queue_reg[1][12]  ( .D(n425), .CPN(Clk_r), .Q(\Queue[1][12] ) );
  FDN1QM1P \Queue_reg[0][12]  ( .D(n457), .CPN(Clk_r), .Q(Packet_Out[12]) );
  FDN1QM1P \Queue_reg[1][11]  ( .D(n424), .CPN(Clk_r), .Q(\Queue[1][11] ) );
  FDN1QM1P \Queue_reg[0][11]  ( .D(n456), .CPN(Clk_r), .Q(Packet_Out[11]) );
  FDN1QM1P \Queue_reg[1][10]  ( .D(n423), .CPN(Clk_r), .Q(\Queue[1][10] ) );
  FDN1QM1P \Queue_reg[0][10]  ( .D(n455), .CPN(Clk_r), .Q(Packet_Out[10]) );
  FDN1QM1P \Queue_reg[1][9]  ( .D(n422), .CPN(Clk_r), .Q(\Queue[1][9] ) );
  FDN1QM1P \Queue_reg[0][9]  ( .D(n454), .CPN(Clk_r), .Q(Packet_Out[9]) );
  FDN1QM1P \Queue_reg[1][8]  ( .D(n421), .CPN(Clk_r), .Q(\Queue[1][8] ) );
  FDN1QM1P \Queue_reg[0][8]  ( .D(n453), .CPN(Clk_r), .Q(Packet_Out[8]) );
  FDN1QM1P \Queue_reg[1][7]  ( .D(n420), .CPN(Clk_r), .Q(\Queue[1][7] ) );
  FDN1QM1P \Queue_reg[0][7]  ( .D(n452), .CPN(Clk_r), .Q(Packet_Out[7]) );
  FDN1QM1P \Queue_reg[1][6]  ( .D(n419), .CPN(Clk_r), .Q(\Queue[1][6] ) );
  FDN1QM1P \Queue_reg[0][6]  ( .D(n451), .CPN(Clk_r), .Q(Packet_Out[6]) );
  FDN1QM1P \Queue_reg[1][5]  ( .D(n418), .CPN(Clk_r), .Q(\Queue[1][5] ) );
  FDN1QM1P \Queue_reg[0][5]  ( .D(n450), .CPN(Clk_r), .Q(Packet_Out[5]) );
  FDN1QM1P \Queue_reg[1][4]  ( .D(n417), .CPN(Clk_r), .Q(\Queue[1][4] ) );
  FDN1QM1P \Queue_reg[0][4]  ( .D(n449), .CPN(Clk_r), .Q(Packet_Out[4]) );
  FDN1QM1P \Queue_reg[1][3]  ( .D(n416), .CPN(Clk_r), .Q(\Queue[1][3] ) );
  FDN1QM1P \Queue_reg[0][3]  ( .D(n448), .CPN(Clk_r), .Q(Packet_Out[3]) );
  FDN1QM1P \Queue_reg[1][2]  ( .D(n415), .CPN(Clk_r), .Q(\Queue[1][2] ) );
  FDN1QM1P \Queue_reg[0][2]  ( .D(n447), .CPN(Clk_r), .Q(Packet_Out[2]) );
  FDN1QM1P \Queue_reg[1][1]  ( .D(n414), .CPN(Clk_r), .Q(\Queue[1][1] ) );
  FDN1QM1P \Queue_reg[0][1]  ( .D(n446), .CPN(Clk_r), .Q(Packet_Out[1]) );
  FDN1QM1P \Queue_reg[1][0]  ( .D(n413), .CPN(Clk_r), .Q(\Queue[1][0] ) );
  FDN1QM1P \Queue_reg[0][0]  ( .D(n445), .CPN(Clk_r), .Q(Packet_Out[0]) );
  FDN2QM1P Empty_reg ( .D(n542), .CPN(Clk_r), .CD(Rst_n), .Q(n541) );
  N1M1P U3 ( .A(Read_Ack), .Z(n137) );
  BUFM2P U4 ( .A(n95), .Z(n3) );
  AOI21M1P U5 ( .A(Write_Ack), .B(n100), .C(n141), .Z(n57) );
  OAI211M4P U6 ( .A(n376), .B(n137), .C(Write_Ack), .D(n62), .Z(n97) );
  OAI211M4P U7 ( .A(n140), .B(n139), .C(Rst_n), .D(n138), .Z(n206) );
  OAI211M4P U8 ( .A(n100), .B(n139), .C(Rst_n), .D(n138), .Z(n133) );
  NR2I1M8P U9 ( .A(n61), .B(n21), .Z(n20) );
  AOI21M2P U10 ( .A(Write_Ack), .B(n142), .C(n141), .Z(n205) );
  AOI21M2P U11 ( .A(Write_Ack), .B(n140), .C(n141), .Z(n132) );
  OAI211M4P U12 ( .A(n100), .B(n137), .C(Write_Ack), .D(n24), .Z(n59) );
  OAI211M4P U13 ( .A(n140), .B(n137), .C(Write_Ack), .D(n98), .Z(n135) );
  OAI211M4P U14 ( .A(n142), .B(n137), .C(Write_Ack), .D(n136), .Z(n208) );
  N1M1P U15 ( .A(Write_Ack), .Z(n99) );
  ND2M1P U16 ( .A(n18), .B(Rst_n), .Z(n61) );
  N1M2P U17 ( .A(n18), .Z(n139) );
  NR2FM1P U18 ( .A(Read_Ack), .B(n99), .Z(n18) );
  NR3M1P U19 ( .A(Count[0]), .B(Count[2]), .C(n22), .Z(n100) );
  NR3M1P U20 ( .A(Count[0]), .B(Count[1]), .C(n19), .Z(n142) );
  NR3M1P U21 ( .A(n23), .B(Count[2]), .C(Count[1]), .Z(n376) );
  NR3M1P U22 ( .A(Count[2]), .B(n23), .C(n22), .Z(n140) );
  N1M1P U23 ( .A(Count[1]), .Z(n22) );
  N1M1P U24 ( .A(Count[0]), .Z(n23) );
  N1M1P U25 ( .A(Count[2]), .Z(n19) );
  BUFM2P U26 ( .A(n132), .Z(n11) );
  BUFM2P U27 ( .A(n205), .Z(n12) );
  ND2M2P U28 ( .A(Read_Ack), .B(Rst_n), .Z(n141) );
  BUFM2P U29 ( .A(n57), .Z(n7) );
  BUFM2P U30 ( .A(n94), .Z(n9) );
  BUFM2P U31 ( .A(n94), .Z(n10) );
  N1M2P U32 ( .A(n62), .Z(n94) );
  BUFM2P U33 ( .A(n56), .Z(n5) );
  BUFM2P U34 ( .A(n56), .Z(n4) );
  BUFM2P U35 ( .A(n56), .Z(n6) );
  BUFM2P U36 ( .A(n57), .Z(n8) );
  NR2M1P U37 ( .A(n137), .B(Write_Ack), .Z(n375) );
  NR2M1P U38 ( .A(n18), .B(n375), .Z(n374) );
  AOI22CDNM1P U39 ( .A(n374), .B(n23), .C(n374), .D(n23), .Z(n377) );
  N1M1P U40 ( .A(n375), .Z(n17) );
  AOI22M1P U41 ( .A(Count[0]), .B(n139), .C(n17), .D(n23), .Z(n14) );
  AOI22CDNM1P U42 ( .A(Count[1]), .B(n14), .C(n14), .D(Count[1]), .Z(n378) );
  ND3M1P U43 ( .A(n23), .B(n19), .C(n22), .Z(n60) );
  ND2M1P U44 ( .A(Count[1]), .B(Read_Ack), .Z(n13) );
  OAI211M1P U45 ( .A(Count[1]), .B(n139), .C(n14), .D(n13), .Z(n15) );
  AOI22M1P U46 ( .A(n18), .B(n140), .C(Count[2]), .D(n15), .Z(n16) );
  OAI21M1P U47 ( .A(n60), .B(n17), .C(n16), .Z(n379) );
  N1M1P U48 ( .A(n142), .Z(n21) );
  N1M1P U49 ( .A(Packet_In[31]), .Z(n373) );
  AOI22CDNM1P U50 ( .A(n20), .B(n373), .C(\Queue[4][31] ), .D(n20), .Z(n380)
         );
  N1M1P U51 ( .A(Packet_In[0]), .Z(n144) );
  AOI22CDNM1P U52 ( .A(n20), .B(n144), .C(\Queue[4][0] ), .D(n20), .Z(n381) );
  N1M1P U53 ( .A(Packet_In[1]), .Z(n146) );
  AOI22CDNM1P U54 ( .A(n20), .B(n146), .C(\Queue[4][1] ), .D(n20), .Z(n382) );
  N1M1P U55 ( .A(Packet_In[2]), .Z(n148) );
  AOI22CDNM1P U56 ( .A(n20), .B(n148), .C(\Queue[4][2] ), .D(n20), .Z(n383) );
  N1M1P U57 ( .A(Packet_In[3]), .Z(n150) );
  AOI22CDNM1P U58 ( .A(n20), .B(n150), .C(\Queue[4][3] ), .D(n20), .Z(n384) );
  N1M1P U59 ( .A(Packet_In[4]), .Z(n152) );
  AOI22CDNM1P U60 ( .A(n20), .B(n152), .C(\Queue[4][4] ), .D(n20), .Z(n385) );
  N1M1P U61 ( .A(Packet_In[5]), .Z(n154) );
  AOI22CDNM1P U62 ( .A(n20), .B(n154), .C(\Queue[4][5] ), .D(n20), .Z(n386) );
  N1M1P U63 ( .A(Packet_In[6]), .Z(n156) );
  AOI22CDNM1P U64 ( .A(n20), .B(n156), .C(\Queue[4][6] ), .D(n20), .Z(n387) );
  N1M1P U65 ( .A(Packet_In[7]), .Z(n158) );
  AOI22CDNM1P U66 ( .A(n20), .B(n158), .C(\Queue[4][7] ), .D(n20), .Z(n388) );
  N1M1P U67 ( .A(Packet_In[8]), .Z(n160) );
  AOI22CDNM1P U68 ( .A(n20), .B(n160), .C(\Queue[4][8] ), .D(n20), .Z(n389) );
  N1M1P U69 ( .A(Packet_In[9]), .Z(n162) );
  AOI22CDNM1P U70 ( .A(n20), .B(n162), .C(\Queue[4][9] ), .D(n20), .Z(n390) );
  N1M1P U71 ( .A(Packet_In[10]), .Z(n164) );
  AOI22CDNM1P U72 ( .A(n20), .B(n164), .C(\Queue[4][10] ), .D(n20), .Z(n391)
         );
  N1M1P U73 ( .A(Packet_In[11]), .Z(n166) );
  AOI22CDNM1P U74 ( .A(n20), .B(n166), .C(\Queue[4][11] ), .D(n20), .Z(n392)
         );
  N1M1P U75 ( .A(Packet_In[12]), .Z(n168) );
  AOI22CDNM1P U76 ( .A(n20), .B(n168), .C(\Queue[4][12] ), .D(n20), .Z(n393)
         );
  N1M1P U77 ( .A(Packet_In[13]), .Z(n170) );
  AOI22CDNM1P U78 ( .A(n20), .B(n170), .C(\Queue[4][13] ), .D(n20), .Z(n394)
         );
  N1M1P U79 ( .A(Packet_In[14]), .Z(n172) );
  AOI22CDNM1P U80 ( .A(n20), .B(n172), .C(\Queue[4][14] ), .D(n20), .Z(n395)
         );
  N1M1P U81 ( .A(Packet_In[15]), .Z(n174) );
  AOI22CDNM1P U82 ( .A(n20), .B(n174), .C(\Queue[4][15] ), .D(n20), .Z(n396)
         );
  N1M1P U83 ( .A(Packet_In[16]), .Z(n176) );
  AOI22CDNM1P U84 ( .A(n20), .B(n176), .C(\Queue[4][16] ), .D(n20), .Z(n397)
         );
  N1M1P U85 ( .A(Packet_In[17]), .Z(n178) );
  AOI22CDNM1P U86 ( .A(n20), .B(n178), .C(\Queue[4][17] ), .D(n20), .Z(n398)
         );
  N1M1P U87 ( .A(Packet_In[18]), .Z(n180) );
  AOI22CDNM1P U88 ( .A(n20), .B(n180), .C(\Queue[4][18] ), .D(n20), .Z(n399)
         );
  N1M1P U89 ( .A(Packet_In[19]), .Z(n182) );
  AOI22CDNM1P U90 ( .A(n20), .B(n182), .C(\Queue[4][19] ), .D(n20), .Z(n400)
         );
  N1M1P U91 ( .A(Packet_In[20]), .Z(n184) );
  AOI22CDNM1P U92 ( .A(n20), .B(n184), .C(\Queue[4][20] ), .D(n20), .Z(n401)
         );
  N1M1P U93 ( .A(Packet_In[21]), .Z(n186) );
  AOI22CDNM1P U94 ( .A(n20), .B(n186), .C(\Queue[4][21] ), .D(n20), .Z(n402)
         );
  N1M1P U95 ( .A(Packet_In[22]), .Z(n188) );
  AOI22CDNM1P U96 ( .A(n20), .B(n188), .C(\Queue[4][22] ), .D(n20), .Z(n403)
         );
  N1M1P U97 ( .A(Packet_In[23]), .Z(n190) );
  AOI22CDNM1P U98 ( .A(n20), .B(n190), .C(\Queue[4][23] ), .D(n20), .Z(n404)
         );
  N1M1P U99 ( .A(Packet_In[24]), .Z(n192) );
  AOI22CDNM1P U100 ( .A(n20), .B(n192), .C(\Queue[4][24] ), .D(n20), .Z(n405)
         );
  N1M1P U101 ( .A(Packet_In[25]), .Z(n194) );
  AOI22CDNM1P U102 ( .A(n20), .B(n194), .C(\Queue[4][25] ), .D(n20), .Z(n406)
         );
  N1M1P U103 ( .A(Packet_In[26]), .Z(n196) );
  AOI22CDNM1P U104 ( .A(n20), .B(n196), .C(\Queue[4][26] ), .D(n20), .Z(n407)
         );
  N1M1P U105 ( .A(Packet_In[27]), .Z(n198) );
  AOI22CDNM1P U106 ( .A(n20), .B(n198), .C(\Queue[4][27] ), .D(n20), .Z(n408)
         );
  N1M1P U107 ( .A(Packet_In[28]), .Z(n200) );
  AOI22CDNM1P U108 ( .A(n20), .B(n200), .C(\Queue[4][28] ), .D(n20), .Z(n409)
         );
  N1M1P U109 ( .A(Packet_In[29]), .Z(n202) );
  AOI22CDNM1P U110 ( .A(n20), .B(n202), .C(\Queue[4][29] ), .D(n20), .Z(n410)
         );
  N1M1P U111 ( .A(Packet_In[30]), .Z(n204) );
  AOI22CDNM1P U112 ( .A(n20), .B(n204), .C(\Queue[4][30] ), .D(n20), .Z(n411)
         );
  OAI22CDNM1P U113 ( .A(n139), .B(n21), .C(n374), .D(Full), .Z(n412) );
  OA21M1P U114 ( .A(n139), .B(n376), .C(Rst_n), .Z(n24) );
  OAI21M1P U115 ( .A(Write_Ack), .B(Read_Ack), .C(n24), .Z(n56) );
  AOI22M1P U116 ( .A(\Queue[2][0] ), .B(n8), .C(\Queue[1][0] ), .D(n4), .Z(n25) );
  OAI21M1P U117 ( .A(n144), .B(n59), .C(n25), .Z(n413) );
  AOI22M1P U118 ( .A(n7), .B(\Queue[2][1] ), .C(\Queue[1][1] ), .D(n4), .Z(n26) );
  OAI21M1P U119 ( .A(n59), .B(n146), .C(n26), .Z(n414) );
  AOI22M1P U120 ( .A(n8), .B(\Queue[2][2] ), .C(\Queue[1][2] ), .D(n4), .Z(n27) );
  OAI21M1P U121 ( .A(n59), .B(n148), .C(n27), .Z(n415) );
  AOI22M1P U122 ( .A(n8), .B(\Queue[2][3] ), .C(\Queue[1][3] ), .D(n4), .Z(n28) );
  OAI21M1P U123 ( .A(n59), .B(n150), .C(n28), .Z(n416) );
  AOI22M1P U124 ( .A(n8), .B(\Queue[2][4] ), .C(\Queue[1][4] ), .D(n4), .Z(n29) );
  OAI21M1P U125 ( .A(n59), .B(n152), .C(n29), .Z(n417) );
  AOI22M1P U126 ( .A(n8), .B(\Queue[2][5] ), .C(\Queue[1][5] ), .D(n4), .Z(n30) );
  OAI21M1P U127 ( .A(n59), .B(n154), .C(n30), .Z(n418) );
  AOI22M1P U128 ( .A(n8), .B(\Queue[2][6] ), .C(\Queue[1][6] ), .D(n4), .Z(n31) );
  OAI21M1P U129 ( .A(n59), .B(n156), .C(n31), .Z(n419) );
  AOI22M1P U130 ( .A(n8), .B(\Queue[2][7] ), .C(\Queue[1][7] ), .D(n4), .Z(n32) );
  OAI21M1P U131 ( .A(n59), .B(n158), .C(n32), .Z(n420) );
  AOI22M1P U132 ( .A(n8), .B(\Queue[2][8] ), .C(\Queue[1][8] ), .D(n4), .Z(n33) );
  OAI21M1P U133 ( .A(n59), .B(n160), .C(n33), .Z(n421) );
  AOI22M1P U134 ( .A(n8), .B(\Queue[2][9] ), .C(\Queue[1][9] ), .D(n5), .Z(n34) );
  OAI21M1P U135 ( .A(n59), .B(n162), .C(n34), .Z(n422) );
  AOI22M1P U136 ( .A(n8), .B(\Queue[2][10] ), .C(\Queue[1][10] ), .D(n5), .Z(
        n35) );
  OAI21M1P U137 ( .A(n59), .B(n164), .C(n35), .Z(n423) );
  AOI22M1P U138 ( .A(n8), .B(\Queue[2][11] ), .C(\Queue[1][11] ), .D(n5), .Z(
        n36) );
  OAI21M1P U139 ( .A(n59), .B(n166), .C(n36), .Z(n424) );
  AOI22M1P U140 ( .A(n7), .B(\Queue[2][12] ), .C(\Queue[1][12] ), .D(n5), .Z(
        n37) );
  OAI21M1P U141 ( .A(n59), .B(n168), .C(n37), .Z(n425) );
  AOI22M1P U142 ( .A(n7), .B(\Queue[2][13] ), .C(\Queue[1][13] ), .D(n5), .Z(
        n38) );
  OAI21M1P U143 ( .A(n59), .B(n170), .C(n38), .Z(n426) );
  AOI22M1P U144 ( .A(n7), .B(\Queue[2][14] ), .C(\Queue[1][14] ), .D(n5), .Z(
        n39) );
  OAI21M1P U145 ( .A(n59), .B(n172), .C(n39), .Z(n427) );
  AOI22M1P U146 ( .A(n7), .B(\Queue[2][15] ), .C(\Queue[1][15] ), .D(n5), .Z(
        n40) );
  OAI21M1P U147 ( .A(n59), .B(n174), .C(n40), .Z(n428) );
  AOI22M1P U148 ( .A(n7), .B(\Queue[2][16] ), .C(\Queue[1][16] ), .D(n5), .Z(
        n41) );
  OAI21M1P U149 ( .A(n59), .B(n176), .C(n41), .Z(n429) );
  AOI22M1P U150 ( .A(n7), .B(\Queue[2][17] ), .C(\Queue[1][17] ), .D(n5), .Z(
        n42) );
  OAI21M1P U151 ( .A(n59), .B(n178), .C(n42), .Z(n430) );
  AOI22M1P U152 ( .A(n7), .B(\Queue[2][18] ), .C(\Queue[1][18] ), .D(n6), .Z(
        n43) );
  OAI21M1P U153 ( .A(n59), .B(n180), .C(n43), .Z(n431) );
  AOI22M1P U154 ( .A(n7), .B(\Queue[2][19] ), .C(\Queue[1][19] ), .D(n6), .Z(
        n44) );
  OAI21M1P U155 ( .A(n59), .B(n182), .C(n44), .Z(n432) );
  AOI22M1P U156 ( .A(n7), .B(\Queue[2][20] ), .C(\Queue[1][20] ), .D(n6), .Z(
        n45) );
  OAI21M1P U157 ( .A(n59), .B(n184), .C(n45), .Z(n433) );
  AOI22M1P U158 ( .A(n7), .B(\Queue[2][21] ), .C(\Queue[1][21] ), .D(n6), .Z(
        n46) );
  OAI21M1P U159 ( .A(n59), .B(n186), .C(n46), .Z(n434) );
  AOI22M1P U160 ( .A(n8), .B(\Queue[2][22] ), .C(\Queue[1][22] ), .D(n6), .Z(
        n47) );
  OAI21M1P U161 ( .A(n59), .B(n188), .C(n47), .Z(n435) );
  AOI22M1P U162 ( .A(n7), .B(\Queue[2][23] ), .C(\Queue[1][23] ), .D(n6), .Z(
        n48) );
  OAI21M1P U163 ( .A(n59), .B(n190), .C(n48), .Z(n436) );
  AOI22M1P U164 ( .A(n8), .B(\Queue[2][24] ), .C(\Queue[1][24] ), .D(n6), .Z(
        n49) );
  OAI21M1P U165 ( .A(n59), .B(n192), .C(n49), .Z(n437) );
  AOI22M1P U166 ( .A(n57), .B(\Queue[2][25] ), .C(\Queue[1][25] ), .D(n6), .Z(
        n50) );
  OAI21M1P U167 ( .A(n59), .B(n194), .C(n50), .Z(n438) );
  AOI22M1P U168 ( .A(n57), .B(\Queue[2][26] ), .C(\Queue[1][26] ), .D(n6), .Z(
        n51) );
  OAI21M1P U169 ( .A(n59), .B(n196), .C(n51), .Z(n439) );
  AOI22M1P U170 ( .A(n57), .B(\Queue[2][27] ), .C(\Queue[1][27] ), .D(n5), .Z(
        n52) );
  OAI21M1P U171 ( .A(n59), .B(n198), .C(n52), .Z(n440) );
  AOI22M1P U172 ( .A(n57), .B(\Queue[2][28] ), .C(\Queue[1][28] ), .D(n6), .Z(
        n53) );
  OAI21M1P U173 ( .A(n59), .B(n200), .C(n53), .Z(n441) );
  AOI22M1P U174 ( .A(n57), .B(\Queue[2][29] ), .C(\Queue[1][29] ), .D(n4), .Z(
        n54) );
  OAI21M1P U175 ( .A(n59), .B(n202), .C(n54), .Z(n442) );
  AOI22M1P U176 ( .A(n57), .B(\Queue[2][30] ), .C(\Queue[1][30] ), .D(n5), .Z(
        n55) );
  OAI21M1P U177 ( .A(n59), .B(n204), .C(n55), .Z(n443) );
  AOI22M1P U178 ( .A(n57), .B(\Queue[2][31] ), .C(\Queue[1][31] ), .D(n6), .Z(
        n58) );
  OAI21M1P U179 ( .A(n59), .B(n373), .C(n58), .Z(n444) );
  OAI21M1P U180 ( .A(n61), .B(n60), .C(n141), .Z(n62) );
  AOI21M1P U181 ( .A(Write_Ack), .B(n376), .C(n141), .Z(n95) );
  AOI22M1P U182 ( .A(\Queue[1][0] ), .B(n3), .C(n94), .D(Packet_Out[0]), .Z(
        n63) );
  OAI21M1P U183 ( .A(n144), .B(n97), .C(n63), .Z(n445) );
  AOI22M1P U184 ( .A(\Queue[1][1] ), .B(n3), .C(n94), .D(Packet_Out[1]), .Z(
        n64) );
  OAI21M1P U185 ( .A(n146), .B(n97), .C(n64), .Z(n446) );
  AOI22M1P U186 ( .A(\Queue[1][2] ), .B(n3), .C(n94), .D(Packet_Out[2]), .Z(
        n65) );
  OAI21M1P U187 ( .A(n148), .B(n97), .C(n65), .Z(n447) );
  AOI22M1P U188 ( .A(\Queue[1][3] ), .B(n3), .C(n94), .D(Packet_Out[3]), .Z(
        n66) );
  OAI21M1P U189 ( .A(n150), .B(n97), .C(n66), .Z(n448) );
  AOI22M1P U190 ( .A(\Queue[1][4] ), .B(n3), .C(n94), .D(Packet_Out[4]), .Z(
        n67) );
  OAI21M1P U191 ( .A(n152), .B(n97), .C(n67), .Z(n449) );
  AOI22M1P U192 ( .A(\Queue[1][5] ), .B(n3), .C(n94), .D(Packet_Out[5]), .Z(
        n68) );
  OAI21M1P U193 ( .A(n154), .B(n97), .C(n68), .Z(n450) );
  AOI22M1P U194 ( .A(\Queue[1][6] ), .B(n3), .C(n94), .D(Packet_Out[6]), .Z(
        n69) );
  OAI21M1P U195 ( .A(n156), .B(n97), .C(n69), .Z(n451) );
  AOI22M1P U196 ( .A(\Queue[1][7] ), .B(n3), .C(n94), .D(Packet_Out[7]), .Z(
        n70) );
  OAI21M1P U197 ( .A(n158), .B(n97), .C(n70), .Z(n452) );
  AOI22M1P U198 ( .A(\Queue[1][8] ), .B(n3), .C(n94), .D(Packet_Out[8]), .Z(
        n71) );
  OAI21M1P U199 ( .A(n160), .B(n97), .C(n71), .Z(n453) );
  AOI22M1P U200 ( .A(\Queue[1][9] ), .B(n3), .C(n94), .D(Packet_Out[9]), .Z(
        n72) );
  OAI21M1P U201 ( .A(n162), .B(n97), .C(n72), .Z(n454) );
  AOI22M1P U202 ( .A(\Queue[1][10] ), .B(n3), .C(n9), .D(Packet_Out[10]), .Z(
        n73) );
  OAI21M1P U203 ( .A(n164), .B(n97), .C(n73), .Z(n455) );
  AOI22M1P U204 ( .A(\Queue[1][11] ), .B(n3), .C(n9), .D(Packet_Out[11]), .Z(
        n74) );
  OAI21M1P U205 ( .A(n166), .B(n97), .C(n74), .Z(n456) );
  AOI22M1P U206 ( .A(\Queue[1][12] ), .B(n3), .C(n9), .D(Packet_Out[12]), .Z(
        n75) );
  OAI21M1P U207 ( .A(n168), .B(n97), .C(n75), .Z(n457) );
  AOI22M1P U208 ( .A(\Queue[1][13] ), .B(n3), .C(n9), .D(Packet_Out[13]), .Z(
        n76) );
  OAI21M1P U209 ( .A(n170), .B(n97), .C(n76), .Z(n458) );
  AOI22M1P U210 ( .A(\Queue[1][14] ), .B(n3), .C(n9), .D(Packet_Out[14]), .Z(
        n77) );
  OAI21M1P U211 ( .A(n172), .B(n97), .C(n77), .Z(n459) );
  AOI22M1P U212 ( .A(\Queue[1][15] ), .B(n3), .C(n9), .D(Packet_Out[15]), .Z(
        n78) );
  OAI21M1P U213 ( .A(n174), .B(n97), .C(n78), .Z(n460) );
  AOI22M1P U214 ( .A(\Queue[1][16] ), .B(n3), .C(n9), .D(Packet_Out[16]), .Z(
        n79) );
  OAI21M1P U215 ( .A(n176), .B(n97), .C(n79), .Z(n461) );
  AOI22M1P U216 ( .A(\Queue[1][17] ), .B(n3), .C(n9), .D(Packet_Out[17]), .Z(
        n80) );
  OAI21M1P U217 ( .A(n178), .B(n97), .C(n80), .Z(n462) );
  AOI22M1P U218 ( .A(\Queue[1][18] ), .B(n3), .C(n9), .D(Packet_Out[18]), .Z(
        n81) );
  OAI21M1P U219 ( .A(n180), .B(n97), .C(n81), .Z(n463) );
  AOI22M1P U220 ( .A(\Queue[1][19] ), .B(n3), .C(n9), .D(Packet_Out[19]), .Z(
        n82) );
  OAI21M1P U221 ( .A(n182), .B(n97), .C(n82), .Z(n464) );
  AOI22M1P U222 ( .A(\Queue[1][20] ), .B(n3), .C(n10), .D(Packet_Out[20]), .Z(
        n83) );
  OAI21M1P U223 ( .A(n184), .B(n97), .C(n83), .Z(n465) );
  AOI22M1P U224 ( .A(\Queue[1][21] ), .B(n3), .C(n10), .D(Packet_Out[21]), .Z(
        n84) );
  OAI21M1P U225 ( .A(n186), .B(n97), .C(n84), .Z(n466) );
  AOI22M1P U226 ( .A(\Queue[1][22] ), .B(n3), .C(n10), .D(Packet_Out[22]), .Z(
        n85) );
  OAI21M1P U227 ( .A(n188), .B(n97), .C(n85), .Z(n467) );
  AOI22M1P U228 ( .A(\Queue[1][23] ), .B(n3), .C(n10), .D(Packet_Out[23]), .Z(
        n86) );
  OAI21M1P U229 ( .A(n190), .B(n97), .C(n86), .Z(n468) );
  AOI22M1P U230 ( .A(\Queue[1][24] ), .B(n3), .C(n10), .D(Packet_Out[24]), .Z(
        n87) );
  OAI21M1P U231 ( .A(n192), .B(n97), .C(n87), .Z(n469) );
  AOI22M1P U232 ( .A(\Queue[1][25] ), .B(n3), .C(n10), .D(Packet_Out[25]), .Z(
        n88) );
  OAI21M1P U233 ( .A(n194), .B(n97), .C(n88), .Z(n470) );
  AOI22M1P U234 ( .A(\Queue[1][26] ), .B(n3), .C(n10), .D(Packet_Out[26]), .Z(
        n89) );
  OAI21M1P U235 ( .A(n196), .B(n97), .C(n89), .Z(n471) );
  AOI22M1P U236 ( .A(\Queue[1][27] ), .B(n3), .C(n10), .D(Packet_Out[27]), .Z(
        n90) );
  OAI21M1P U237 ( .A(n198), .B(n97), .C(n90), .Z(n472) );
  AOI22M1P U238 ( .A(\Queue[1][28] ), .B(n3), .C(n10), .D(Packet_Out[28]), .Z(
        n91) );
  OAI21M1P U239 ( .A(n200), .B(n97), .C(n91), .Z(n473) );
  AOI22M1P U240 ( .A(\Queue[1][29] ), .B(n3), .C(n10), .D(Packet_Out[29]), .Z(
        n92) );
  OAI21M1P U241 ( .A(n202), .B(n97), .C(n92), .Z(n474) );
  AOI22M1P U242 ( .A(\Queue[1][30] ), .B(n95), .C(n9), .D(Packet_Out[30]), .Z(
        n93) );
  OAI21M1P U243 ( .A(n204), .B(n97), .C(n93), .Z(n475) );
  AOI22M1P U244 ( .A(\Queue[1][31] ), .B(n95), .C(n10), .D(Packet_Out[31]), 
        .Z(n96) );
  OAI21M1P U245 ( .A(n373), .B(n97), .C(n96), .Z(n476) );
  OA21M1P U246 ( .A(n139), .B(n100), .C(Rst_n), .Z(n98) );
  ND2M1P U247 ( .A(n99), .B(n137), .Z(n138) );
  AOI22M1P U248 ( .A(\Queue[2][0] ), .B(n133), .C(\Queue[3][0] ), .D(n11), .Z(
        n101) );
  OAI21M1P U249 ( .A(n144), .B(n135), .C(n101), .Z(n477) );
  AOI22M1P U250 ( .A(\Queue[2][1] ), .B(n133), .C(n132), .D(\Queue[3][1] ), 
        .Z(n102) );
  OAI21M1P U251 ( .A(n146), .B(n135), .C(n102), .Z(n478) );
  AOI22M1P U252 ( .A(\Queue[2][2] ), .B(n133), .C(n11), .D(\Queue[3][2] ), .Z(
        n103) );
  OAI21M1P U253 ( .A(n148), .B(n135), .C(n103), .Z(n479) );
  AOI22M1P U254 ( .A(\Queue[2][3] ), .B(n133), .C(n11), .D(\Queue[3][3] ), .Z(
        n104) );
  OAI21M1P U255 ( .A(n150), .B(n135), .C(n104), .Z(n480) );
  AOI22M1P U256 ( .A(\Queue[2][4] ), .B(n133), .C(n11), .D(\Queue[3][4] ), .Z(
        n105) );
  OAI21M1P U257 ( .A(n152), .B(n135), .C(n105), .Z(n481) );
  AOI22M1P U258 ( .A(\Queue[2][5] ), .B(n133), .C(n11), .D(\Queue[3][5] ), .Z(
        n106) );
  OAI21M1P U259 ( .A(n154), .B(n135), .C(n106), .Z(n482) );
  AOI22M1P U260 ( .A(\Queue[2][6] ), .B(n133), .C(n11), .D(\Queue[3][6] ), .Z(
        n107) );
  OAI21M1P U261 ( .A(n156), .B(n135), .C(n107), .Z(n483) );
  AOI22M1P U262 ( .A(\Queue[2][7] ), .B(n133), .C(n11), .D(\Queue[3][7] ), .Z(
        n108) );
  OAI21M1P U263 ( .A(n158), .B(n135), .C(n108), .Z(n484) );
  AOI22M1P U264 ( .A(\Queue[2][8] ), .B(n133), .C(n11), .D(\Queue[3][8] ), .Z(
        n109) );
  OAI21M1P U265 ( .A(n160), .B(n135), .C(n109), .Z(n485) );
  AOI22M1P U266 ( .A(\Queue[2][9] ), .B(n133), .C(n11), .D(\Queue[3][9] ), .Z(
        n110) );
  OAI21M1P U267 ( .A(n162), .B(n135), .C(n110), .Z(n486) );
  AOI22M1P U268 ( .A(\Queue[2][10] ), .B(n133), .C(n11), .D(\Queue[3][10] ), 
        .Z(n111) );
  OAI21M1P U269 ( .A(n164), .B(n135), .C(n111), .Z(n487) );
  AOI22M1P U270 ( .A(\Queue[2][11] ), .B(n133), .C(n11), .D(\Queue[3][11] ), 
        .Z(n112) );
  OAI21M1P U271 ( .A(n166), .B(n135), .C(n112), .Z(n488) );
  AOI22M1P U272 ( .A(\Queue[2][12] ), .B(n133), .C(n132), .D(\Queue[3][12] ), 
        .Z(n113) );
  OAI21M1P U273 ( .A(n168), .B(n135), .C(n113), .Z(n489) );
  AOI22M1P U274 ( .A(\Queue[2][13] ), .B(n133), .C(n132), .D(\Queue[3][13] ), 
        .Z(n114) );
  OAI21M1P U275 ( .A(n170), .B(n135), .C(n114), .Z(n490) );
  AOI22M1P U276 ( .A(\Queue[2][14] ), .B(n133), .C(n132), .D(\Queue[3][14] ), 
        .Z(n115) );
  OAI21M1P U277 ( .A(n172), .B(n135), .C(n115), .Z(n491) );
  AOI22M1P U278 ( .A(\Queue[2][15] ), .B(n133), .C(n132), .D(\Queue[3][15] ), 
        .Z(n116) );
  OAI21M1P U279 ( .A(n174), .B(n135), .C(n116), .Z(n492) );
  AOI22M1P U280 ( .A(\Queue[2][16] ), .B(n133), .C(n132), .D(\Queue[3][16] ), 
        .Z(n117) );
  OAI21M1P U281 ( .A(n176), .B(n135), .C(n117), .Z(n493) );
  AOI22M1P U282 ( .A(\Queue[2][17] ), .B(n133), .C(n11), .D(\Queue[3][17] ), 
        .Z(n118) );
  OAI21M1P U283 ( .A(n178), .B(n135), .C(n118), .Z(n494) );
  AOI22M1P U284 ( .A(\Queue[2][18] ), .B(n133), .C(n132), .D(\Queue[3][18] ), 
        .Z(n119) );
  OAI21M1P U285 ( .A(n180), .B(n135), .C(n119), .Z(n495) );
  AOI22M1P U286 ( .A(\Queue[2][19] ), .B(n133), .C(n132), .D(\Queue[3][19] ), 
        .Z(n120) );
  OAI21M1P U287 ( .A(n182), .B(n135), .C(n120), .Z(n496) );
  AOI22M1P U288 ( .A(\Queue[2][20] ), .B(n133), .C(n132), .D(\Queue[3][20] ), 
        .Z(n121) );
  OAI21M1P U289 ( .A(n184), .B(n135), .C(n121), .Z(n497) );
  AOI22M1P U290 ( .A(\Queue[2][21] ), .B(n133), .C(n132), .D(\Queue[3][21] ), 
        .Z(n122) );
  OAI21M1P U291 ( .A(n186), .B(n135), .C(n122), .Z(n498) );
  AOI22M1P U292 ( .A(\Queue[2][22] ), .B(n133), .C(n11), .D(\Queue[3][22] ), 
        .Z(n123) );
  OAI21M1P U293 ( .A(n188), .B(n135), .C(n123), .Z(n499) );
  AOI22M1P U294 ( .A(\Queue[2][23] ), .B(n133), .C(n11), .D(\Queue[3][23] ), 
        .Z(n124) );
  OAI21M1P U295 ( .A(n190), .B(n135), .C(n124), .Z(n500) );
  AOI22M1P U296 ( .A(\Queue[2][24] ), .B(n133), .C(n11), .D(\Queue[3][24] ), 
        .Z(n125) );
  OAI21M1P U297 ( .A(n192), .B(n135), .C(n125), .Z(n501) );
  AOI22M1P U298 ( .A(\Queue[2][25] ), .B(n133), .C(n11), .D(\Queue[3][25] ), 
        .Z(n126) );
  OAI21M1P U299 ( .A(n194), .B(n135), .C(n126), .Z(n502) );
  AOI22M1P U300 ( .A(\Queue[2][26] ), .B(n133), .C(n11), .D(\Queue[3][26] ), 
        .Z(n127) );
  OAI21M1P U301 ( .A(n196), .B(n135), .C(n127), .Z(n503) );
  AOI22M1P U302 ( .A(\Queue[2][27] ), .B(n133), .C(n11), .D(\Queue[3][27] ), 
        .Z(n128) );
  OAI21M1P U303 ( .A(n198), .B(n135), .C(n128), .Z(n504) );
  AOI22M1P U304 ( .A(\Queue[2][28] ), .B(n133), .C(n11), .D(\Queue[3][28] ), 
        .Z(n129) );
  OAI21M1P U305 ( .A(n200), .B(n135), .C(n129), .Z(n505) );
  AOI22M1P U306 ( .A(\Queue[2][29] ), .B(n133), .C(n11), .D(\Queue[3][29] ), 
        .Z(n130) );
  OAI21M1P U307 ( .A(n202), .B(n135), .C(n130), .Z(n506) );
  AOI22M1P U308 ( .A(\Queue[2][30] ), .B(n133), .C(n132), .D(\Queue[3][30] ), 
        .Z(n131) );
  OAI21M1P U309 ( .A(n204), .B(n135), .C(n131), .Z(n507) );
  AOI22M1P U310 ( .A(\Queue[2][31] ), .B(n133), .C(n132), .D(\Queue[3][31] ), 
        .Z(n134) );
  OAI21M1P U311 ( .A(n373), .B(n135), .C(n134), .Z(n508) );
  OA21M1P U312 ( .A(n139), .B(n140), .C(Rst_n), .Z(n136) );
  AOI22M1P U313 ( .A(\Queue[3][0] ), .B(n206), .C(n12), .D(\Queue[4][0] ), .Z(
        n143) );
  OAI21M1P U314 ( .A(n144), .B(n208), .C(n143), .Z(n509) );
  AOI22M1P U315 ( .A(\Queue[3][1] ), .B(n206), .C(n12), .D(\Queue[4][1] ), .Z(
        n145) );
  OAI21M1P U316 ( .A(n146), .B(n208), .C(n145), .Z(n510) );
  AOI22M1P U317 ( .A(\Queue[3][2] ), .B(n206), .C(n12), .D(\Queue[4][2] ), .Z(
        n147) );
  OAI21M1P U318 ( .A(n148), .B(n208), .C(n147), .Z(n511) );
  AOI22M1P U319 ( .A(\Queue[3][3] ), .B(n206), .C(n12), .D(\Queue[4][3] ), .Z(
        n149) );
  OAI21M1P U320 ( .A(n150), .B(n208), .C(n149), .Z(n512) );
  AOI22M1P U321 ( .A(\Queue[3][4] ), .B(n206), .C(n12), .D(\Queue[4][4] ), .Z(
        n151) );
  OAI21M1P U322 ( .A(n152), .B(n208), .C(n151), .Z(n513) );
  AOI22M1P U323 ( .A(\Queue[3][5] ), .B(n206), .C(n12), .D(\Queue[4][5] ), .Z(
        n153) );
  OAI21M1P U324 ( .A(n154), .B(n208), .C(n153), .Z(n514) );
  AOI22M1P U325 ( .A(\Queue[3][6] ), .B(n206), .C(n12), .D(\Queue[4][6] ), .Z(
        n155) );
  OAI21M1P U326 ( .A(n156), .B(n208), .C(n155), .Z(n515) );
  AOI22M1P U327 ( .A(\Queue[3][7] ), .B(n206), .C(n12), .D(\Queue[4][7] ), .Z(
        n157) );
  OAI21M1P U328 ( .A(n158), .B(n208), .C(n157), .Z(n516) );
  AOI22M1P U329 ( .A(\Queue[3][8] ), .B(n206), .C(n205), .D(\Queue[4][8] ), 
        .Z(n159) );
  OAI21M1P U330 ( .A(n160), .B(n208), .C(n159), .Z(n517) );
  AOI22M1P U331 ( .A(\Queue[3][9] ), .B(n206), .C(n205), .D(\Queue[4][9] ), 
        .Z(n161) );
  OAI21M1P U332 ( .A(n162), .B(n208), .C(n161), .Z(n518) );
  AOI22M1P U333 ( .A(\Queue[3][10] ), .B(n206), .C(n12), .D(\Queue[4][10] ), 
        .Z(n163) );
  OAI21M1P U334 ( .A(n164), .B(n208), .C(n163), .Z(n519) );
  AOI22M1P U335 ( .A(\Queue[3][11] ), .B(n206), .C(n205), .D(\Queue[4][11] ), 
        .Z(n165) );
  OAI21M1P U336 ( .A(n166), .B(n208), .C(n165), .Z(n520) );
  AOI22M1P U337 ( .A(\Queue[3][12] ), .B(n206), .C(n12), .D(\Queue[4][12] ), 
        .Z(n167) );
  OAI21M1P U338 ( .A(n168), .B(n208), .C(n167), .Z(n521) );
  AOI22M1P U339 ( .A(\Queue[3][13] ), .B(n206), .C(n12), .D(\Queue[4][13] ), 
        .Z(n169) );
  OAI21M1P U340 ( .A(n170), .B(n208), .C(n169), .Z(n522) );
  AOI22M1P U341 ( .A(\Queue[3][14] ), .B(n206), .C(n12), .D(\Queue[4][14] ), 
        .Z(n171) );
  OAI21M1P U342 ( .A(n172), .B(n208), .C(n171), .Z(n523) );
  AOI22M1P U343 ( .A(\Queue[3][15] ), .B(n206), .C(n12), .D(\Queue[4][15] ), 
        .Z(n173) );
  OAI21M1P U344 ( .A(n174), .B(n208), .C(n173), .Z(n524) );
  AOI22M1P U345 ( .A(\Queue[3][16] ), .B(n206), .C(n12), .D(\Queue[4][16] ), 
        .Z(n175) );
  OAI21M1P U346 ( .A(n176), .B(n208), .C(n175), .Z(n525) );
  AOI22M1P U347 ( .A(\Queue[3][17] ), .B(n206), .C(n12), .D(\Queue[4][17] ), 
        .Z(n177) );
  OAI21M1P U348 ( .A(n178), .B(n208), .C(n177), .Z(n526) );
  AOI22M1P U349 ( .A(\Queue[3][18] ), .B(n206), .C(n12), .D(\Queue[4][18] ), 
        .Z(n179) );
  OAI21M1P U350 ( .A(n180), .B(n208), .C(n179), .Z(n527) );
  AOI22M1P U351 ( .A(\Queue[3][19] ), .B(n206), .C(n12), .D(\Queue[4][19] ), 
        .Z(n181) );
  OAI21M1P U352 ( .A(n182), .B(n208), .C(n181), .Z(n528) );
  AOI22M1P U353 ( .A(\Queue[3][20] ), .B(n206), .C(n205), .D(\Queue[4][20] ), 
        .Z(n183) );
  OAI21M1P U354 ( .A(n184), .B(n208), .C(n183), .Z(n529) );
  AOI22M1P U355 ( .A(\Queue[3][21] ), .B(n206), .C(n205), .D(\Queue[4][21] ), 
        .Z(n185) );
  OAI21M1P U356 ( .A(n186), .B(n208), .C(n185), .Z(n530) );
  AOI22M1P U357 ( .A(\Queue[3][22] ), .B(n206), .C(n205), .D(\Queue[4][22] ), 
        .Z(n187) );
  OAI21M1P U358 ( .A(n188), .B(n208), .C(n187), .Z(n531) );
  AOI22M1P U359 ( .A(\Queue[3][23] ), .B(n206), .C(n205), .D(\Queue[4][23] ), 
        .Z(n189) );
  OAI21M1P U360 ( .A(n190), .B(n208), .C(n189), .Z(n532) );
  AOI22M1P U361 ( .A(\Queue[3][24] ), .B(n206), .C(n205), .D(\Queue[4][24] ), 
        .Z(n191) );
  OAI21M1P U362 ( .A(n192), .B(n208), .C(n191), .Z(n533) );
  AOI22M1P U363 ( .A(\Queue[3][25] ), .B(n206), .C(n205), .D(\Queue[4][25] ), 
        .Z(n193) );
  OAI21M1P U364 ( .A(n194), .B(n208), .C(n193), .Z(n534) );
  AOI22M1P U365 ( .A(\Queue[3][26] ), .B(n206), .C(n205), .D(\Queue[4][26] ), 
        .Z(n195) );
  OAI21M1P U366 ( .A(n196), .B(n208), .C(n195), .Z(n535) );
  AOI22M1P U367 ( .A(\Queue[3][27] ), .B(n206), .C(n205), .D(\Queue[4][27] ), 
        .Z(n197) );
  OAI21M1P U368 ( .A(n198), .B(n208), .C(n197), .Z(n536) );
  AOI22M1P U369 ( .A(\Queue[3][28] ), .B(n206), .C(n12), .D(\Queue[4][28] ), 
        .Z(n199) );
  OAI21M1P U370 ( .A(n200), .B(n208), .C(n199), .Z(n537) );
  AOI22M1P U371 ( .A(\Queue[3][29] ), .B(n206), .C(n205), .D(\Queue[4][29] ), 
        .Z(n201) );
  OAI21M1P U372 ( .A(n202), .B(n208), .C(n201), .Z(n538) );
  AOI22M1P U373 ( .A(\Queue[3][30] ), .B(n206), .C(n12), .D(\Queue[4][30] ), 
        .Z(n203) );
  OAI21M1P U374 ( .A(n204), .B(n208), .C(n203), .Z(n539) );
  AOI22M1P U375 ( .A(\Queue[3][31] ), .B(n206), .C(n12), .D(\Queue[4][31] ), 
        .Z(n207) );
  OAI21M1P U376 ( .A(n373), .B(n208), .C(n207), .Z(n540) );
  N1M1P U377 ( .A(n541), .Z(Empty) );
  AOI22M1P U378 ( .A(n376), .B(n375), .C(n374), .D(Empty), .Z(n542) );
endmodule


module Packet_Queue_4 ( Clk_r, Rst_n, Packet_In, Read_Ack, Write_Ack, 
        Packet_Out, Empty, Full );
  input [31:0] Packet_In;
  output [31:0] Packet_Out;
  input Clk_r, Rst_n, Read_Ack, Write_Ack;
  output Empty, Full;
  wire   \Queue[4][31] , \Queue[4][30] , \Queue[4][29] , \Queue[4][28] ,
         \Queue[4][27] , \Queue[4][26] , \Queue[4][25] , \Queue[4][24] ,
         \Queue[4][23] , \Queue[4][22] , \Queue[4][21] , \Queue[4][20] ,
         \Queue[4][19] , \Queue[4][18] , \Queue[4][17] , \Queue[4][16] ,
         \Queue[4][15] , \Queue[4][14] , \Queue[4][13] , \Queue[4][12] ,
         \Queue[4][11] , \Queue[4][10] , \Queue[4][9] , \Queue[4][8] ,
         \Queue[4][7] , \Queue[4][6] , \Queue[4][5] , \Queue[4][4] ,
         \Queue[4][3] , \Queue[4][2] , \Queue[4][1] , \Queue[4][0] ,
         \Queue[3][31] , \Queue[3][30] , \Queue[3][29] , \Queue[3][28] ,
         \Queue[3][27] , \Queue[3][26] , \Queue[3][25] , \Queue[3][24] ,
         \Queue[3][23] , \Queue[3][22] , \Queue[3][21] , \Queue[3][20] ,
         \Queue[3][19] , \Queue[3][18] , \Queue[3][17] , \Queue[3][16] ,
         \Queue[3][15] , \Queue[3][14] , \Queue[3][13] , \Queue[3][12] ,
         \Queue[3][11] , \Queue[3][10] , \Queue[3][9] , \Queue[3][8] ,
         \Queue[3][7] , \Queue[3][6] , \Queue[3][5] , \Queue[3][4] ,
         \Queue[3][3] , \Queue[3][2] , \Queue[3][1] , \Queue[3][0] ,
         \Queue[2][31] , \Queue[2][30] , \Queue[2][29] , \Queue[2][28] ,
         \Queue[2][27] , \Queue[2][26] , \Queue[2][25] , \Queue[2][24] ,
         \Queue[2][23] , \Queue[2][22] , \Queue[2][21] , \Queue[2][20] ,
         \Queue[2][19] , \Queue[2][18] , \Queue[2][17] , \Queue[2][16] ,
         \Queue[2][15] , \Queue[2][14] , \Queue[2][13] , \Queue[2][12] ,
         \Queue[2][11] , \Queue[2][10] , \Queue[2][9] , \Queue[2][8] ,
         \Queue[2][7] , \Queue[2][6] , \Queue[2][5] , \Queue[2][4] ,
         \Queue[2][3] , \Queue[2][2] , \Queue[2][1] , \Queue[2][0] ,
         \Queue[1][31] , \Queue[1][30] , \Queue[1][29] , \Queue[1][28] ,
         \Queue[1][27] , \Queue[1][26] , \Queue[1][25] , \Queue[1][24] ,
         \Queue[1][23] , \Queue[1][22] , \Queue[1][21] , \Queue[1][20] ,
         \Queue[1][19] , \Queue[1][18] , \Queue[1][17] , \Queue[1][16] ,
         \Queue[1][15] , \Queue[1][14] , \Queue[1][13] , \Queue[1][12] ,
         \Queue[1][11] , \Queue[1][10] , \Queue[1][9] , \Queue[1][8] ,
         \Queue[1][7] , \Queue[1][6] , \Queue[1][5] , \Queue[1][4] ,
         \Queue[1][3] , \Queue[1][2] , \Queue[1][1] , \Queue[1][0] , n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550;
  wire   [2:0] Count;

  FDN2QM1P \Count_reg[0]  ( .D(n385), .CPN(Clk_r), .CD(Rst_n), .Q(Count[0]) );
  FDN2QM1P \Count_reg[1]  ( .D(n386), .CPN(Clk_r), .CD(Rst_n), .Q(Count[1]) );
  FDN2QM1P \Count_reg[2]  ( .D(n387), .CPN(Clk_r), .CD(Rst_n), .Q(Count[2]) );
  FDN1QM1P \Queue_reg[4][30]  ( .D(n419), .CPN(Clk_r), .Q(\Queue[4][30] ) );
  FDN1QM1P \Queue_reg[3][30]  ( .D(n547), .CPN(Clk_r), .Q(\Queue[3][30] ) );
  FDN1QM1P \Queue_reg[2][30]  ( .D(n515), .CPN(Clk_r), .Q(\Queue[2][30] ) );
  FDN1QM1P \Queue_reg[4][29]  ( .D(n418), .CPN(Clk_r), .Q(\Queue[4][29] ) );
  FDN1QM1P \Queue_reg[3][29]  ( .D(n546), .CPN(Clk_r), .Q(\Queue[3][29] ) );
  FDN1QM1P \Queue_reg[2][29]  ( .D(n514), .CPN(Clk_r), .Q(\Queue[2][29] ) );
  FDN1QM1P \Queue_reg[4][28]  ( .D(n417), .CPN(Clk_r), .Q(\Queue[4][28] ) );
  FDN1QM1P \Queue_reg[3][28]  ( .D(n545), .CPN(Clk_r), .Q(\Queue[3][28] ) );
  FDN1QM1P \Queue_reg[2][28]  ( .D(n513), .CPN(Clk_r), .Q(\Queue[2][28] ) );
  FDN1QM1P \Queue_reg[4][27]  ( .D(n416), .CPN(Clk_r), .Q(\Queue[4][27] ) );
  FDN1QM1P \Queue_reg[3][27]  ( .D(n544), .CPN(Clk_r), .Q(\Queue[3][27] ) );
  FDN1QM1P \Queue_reg[2][27]  ( .D(n512), .CPN(Clk_r), .Q(\Queue[2][27] ) );
  FDN1QM1P \Queue_reg[4][26]  ( .D(n415), .CPN(Clk_r), .Q(\Queue[4][26] ) );
  FDN1QM1P \Queue_reg[3][26]  ( .D(n543), .CPN(Clk_r), .Q(\Queue[3][26] ) );
  FDN1QM1P \Queue_reg[2][26]  ( .D(n511), .CPN(Clk_r), .Q(\Queue[2][26] ) );
  FDN1QM1P \Queue_reg[4][25]  ( .D(n414), .CPN(Clk_r), .Q(\Queue[4][25] ) );
  FDN1QM1P \Queue_reg[3][25]  ( .D(n542), .CPN(Clk_r), .Q(\Queue[3][25] ) );
  FDN1QM1P \Queue_reg[2][25]  ( .D(n510), .CPN(Clk_r), .Q(\Queue[2][25] ) );
  FDN1QM1P \Queue_reg[4][24]  ( .D(n413), .CPN(Clk_r), .Q(\Queue[4][24] ) );
  FDN1QM1P \Queue_reg[3][24]  ( .D(n541), .CPN(Clk_r), .Q(\Queue[3][24] ) );
  FDN1QM1P \Queue_reg[2][24]  ( .D(n509), .CPN(Clk_r), .Q(\Queue[2][24] ) );
  FDN1QM1P \Queue_reg[4][23]  ( .D(n412), .CPN(Clk_r), .Q(\Queue[4][23] ) );
  FDN1QM1P \Queue_reg[3][23]  ( .D(n540), .CPN(Clk_r), .Q(\Queue[3][23] ) );
  FDN1QM1P \Queue_reg[2][23]  ( .D(n508), .CPN(Clk_r), .Q(\Queue[2][23] ) );
  FDN1QM1P \Queue_reg[4][22]  ( .D(n411), .CPN(Clk_r), .Q(\Queue[4][22] ) );
  FDN1QM1P \Queue_reg[3][22]  ( .D(n539), .CPN(Clk_r), .Q(\Queue[3][22] ) );
  FDN1QM1P \Queue_reg[2][22]  ( .D(n507), .CPN(Clk_r), .Q(\Queue[2][22] ) );
  FDN1QM1P \Queue_reg[4][21]  ( .D(n410), .CPN(Clk_r), .Q(\Queue[4][21] ) );
  FDN1QM1P \Queue_reg[3][21]  ( .D(n538), .CPN(Clk_r), .Q(\Queue[3][21] ) );
  FDN1QM1P \Queue_reg[2][21]  ( .D(n506), .CPN(Clk_r), .Q(\Queue[2][21] ) );
  FDN1QM1P \Queue_reg[4][20]  ( .D(n409), .CPN(Clk_r), .Q(\Queue[4][20] ) );
  FDN1QM1P \Queue_reg[3][20]  ( .D(n537), .CPN(Clk_r), .Q(\Queue[3][20] ) );
  FDN1QM1P \Queue_reg[2][20]  ( .D(n505), .CPN(Clk_r), .Q(\Queue[2][20] ) );
  FDN1QM1P \Queue_reg[4][19]  ( .D(n408), .CPN(Clk_r), .Q(\Queue[4][19] ) );
  FDN1QM1P \Queue_reg[3][19]  ( .D(n536), .CPN(Clk_r), .Q(\Queue[3][19] ) );
  FDN1QM1P \Queue_reg[2][19]  ( .D(n504), .CPN(Clk_r), .Q(\Queue[2][19] ) );
  FDN1QM1P \Queue_reg[4][18]  ( .D(n407), .CPN(Clk_r), .Q(\Queue[4][18] ) );
  FDN1QM1P \Queue_reg[3][18]  ( .D(n535), .CPN(Clk_r), .Q(\Queue[3][18] ) );
  FDN1QM1P \Queue_reg[2][18]  ( .D(n503), .CPN(Clk_r), .Q(\Queue[2][18] ) );
  FDN1QM1P \Queue_reg[4][17]  ( .D(n406), .CPN(Clk_r), .Q(\Queue[4][17] ) );
  FDN1QM1P \Queue_reg[3][17]  ( .D(n534), .CPN(Clk_r), .Q(\Queue[3][17] ) );
  FDN1QM1P \Queue_reg[2][17]  ( .D(n502), .CPN(Clk_r), .Q(\Queue[2][17] ) );
  FDN1QM1P \Queue_reg[4][16]  ( .D(n405), .CPN(Clk_r), .Q(\Queue[4][16] ) );
  FDN1QM1P \Queue_reg[3][16]  ( .D(n533), .CPN(Clk_r), .Q(\Queue[3][16] ) );
  FDN1QM1P \Queue_reg[2][16]  ( .D(n501), .CPN(Clk_r), .Q(\Queue[2][16] ) );
  FDN1QM1P \Queue_reg[4][15]  ( .D(n404), .CPN(Clk_r), .Q(\Queue[4][15] ) );
  FDN1QM1P \Queue_reg[3][15]  ( .D(n532), .CPN(Clk_r), .Q(\Queue[3][15] ) );
  FDN1QM1P \Queue_reg[2][15]  ( .D(n500), .CPN(Clk_r), .Q(\Queue[2][15] ) );
  FDN1QM1P \Queue_reg[4][14]  ( .D(n403), .CPN(Clk_r), .Q(\Queue[4][14] ) );
  FDN1QM1P \Queue_reg[3][14]  ( .D(n531), .CPN(Clk_r), .Q(\Queue[3][14] ) );
  FDN1QM1P \Queue_reg[2][14]  ( .D(n499), .CPN(Clk_r), .Q(\Queue[2][14] ) );
  FDN1QM1P \Queue_reg[4][13]  ( .D(n402), .CPN(Clk_r), .Q(\Queue[4][13] ) );
  FDN1QM1P \Queue_reg[3][13]  ( .D(n530), .CPN(Clk_r), .Q(\Queue[3][13] ) );
  FDN1QM1P \Queue_reg[2][13]  ( .D(n498), .CPN(Clk_r), .Q(\Queue[2][13] ) );
  FDN1QM1P \Queue_reg[4][12]  ( .D(n401), .CPN(Clk_r), .Q(\Queue[4][12] ) );
  FDN1QM1P \Queue_reg[3][12]  ( .D(n529), .CPN(Clk_r), .Q(\Queue[3][12] ) );
  FDN1QM1P \Queue_reg[2][12]  ( .D(n497), .CPN(Clk_r), .Q(\Queue[2][12] ) );
  FDN1QM1P \Queue_reg[4][11]  ( .D(n400), .CPN(Clk_r), .Q(\Queue[4][11] ) );
  FDN1QM1P \Queue_reg[3][11]  ( .D(n528), .CPN(Clk_r), .Q(\Queue[3][11] ) );
  FDN1QM1P \Queue_reg[2][11]  ( .D(n496), .CPN(Clk_r), .Q(\Queue[2][11] ) );
  FDN1QM1P \Queue_reg[4][10]  ( .D(n399), .CPN(Clk_r), .Q(\Queue[4][10] ) );
  FDN1QM1P \Queue_reg[3][10]  ( .D(n527), .CPN(Clk_r), .Q(\Queue[3][10] ) );
  FDN1QM1P \Queue_reg[2][10]  ( .D(n495), .CPN(Clk_r), .Q(\Queue[2][10] ) );
  FDN1QM1P \Queue_reg[4][9]  ( .D(n398), .CPN(Clk_r), .Q(\Queue[4][9] ) );
  FDN1QM1P \Queue_reg[3][9]  ( .D(n526), .CPN(Clk_r), .Q(\Queue[3][9] ) );
  FDN1QM1P \Queue_reg[2][9]  ( .D(n494), .CPN(Clk_r), .Q(\Queue[2][9] ) );
  FDN1QM1P \Queue_reg[4][8]  ( .D(n397), .CPN(Clk_r), .Q(\Queue[4][8] ) );
  FDN1QM1P \Queue_reg[3][8]  ( .D(n525), .CPN(Clk_r), .Q(\Queue[3][8] ) );
  FDN1QM1P \Queue_reg[2][8]  ( .D(n493), .CPN(Clk_r), .Q(\Queue[2][8] ) );
  FDN1QM1P \Queue_reg[4][7]  ( .D(n396), .CPN(Clk_r), .Q(\Queue[4][7] ) );
  FDN1QM1P \Queue_reg[3][7]  ( .D(n524), .CPN(Clk_r), .Q(\Queue[3][7] ) );
  FDN1QM1P \Queue_reg[2][7]  ( .D(n492), .CPN(Clk_r), .Q(\Queue[2][7] ) );
  FDN1QM1P \Queue_reg[4][6]  ( .D(n395), .CPN(Clk_r), .Q(\Queue[4][6] ) );
  FDN1QM1P \Queue_reg[3][6]  ( .D(n523), .CPN(Clk_r), .Q(\Queue[3][6] ) );
  FDN1QM1P \Queue_reg[2][6]  ( .D(n491), .CPN(Clk_r), .Q(\Queue[2][6] ) );
  FDN1QM1P \Queue_reg[4][5]  ( .D(n394), .CPN(Clk_r), .Q(\Queue[4][5] ) );
  FDN1QM1P \Queue_reg[3][5]  ( .D(n522), .CPN(Clk_r), .Q(\Queue[3][5] ) );
  FDN1QM1P \Queue_reg[2][5]  ( .D(n490), .CPN(Clk_r), .Q(\Queue[2][5] ) );
  FDN1QM1P \Queue_reg[4][4]  ( .D(n393), .CPN(Clk_r), .Q(\Queue[4][4] ) );
  FDN1QM1P \Queue_reg[3][4]  ( .D(n521), .CPN(Clk_r), .Q(\Queue[3][4] ) );
  FDN1QM1P \Queue_reg[2][4]  ( .D(n489), .CPN(Clk_r), .Q(\Queue[2][4] ) );
  FDN1QM1P \Queue_reg[4][3]  ( .D(n392), .CPN(Clk_r), .Q(\Queue[4][3] ) );
  FDN1QM1P \Queue_reg[3][3]  ( .D(n520), .CPN(Clk_r), .Q(\Queue[3][3] ) );
  FDN1QM1P \Queue_reg[2][3]  ( .D(n488), .CPN(Clk_r), .Q(\Queue[2][3] ) );
  FDN1QM1P \Queue_reg[4][2]  ( .D(n391), .CPN(Clk_r), .Q(\Queue[4][2] ) );
  FDN1QM1P \Queue_reg[3][2]  ( .D(n519), .CPN(Clk_r), .Q(\Queue[3][2] ) );
  FDN1QM1P \Queue_reg[2][2]  ( .D(n487), .CPN(Clk_r), .Q(\Queue[2][2] ) );
  FDN1QM1P \Queue_reg[4][1]  ( .D(n390), .CPN(Clk_r), .Q(\Queue[4][1] ) );
  FDN1QM1P \Queue_reg[3][1]  ( .D(n518), .CPN(Clk_r), .Q(\Queue[3][1] ) );
  FDN1QM1P \Queue_reg[2][1]  ( .D(n486), .CPN(Clk_r), .Q(\Queue[2][1] ) );
  FDN1QM1P \Queue_reg[4][0]  ( .D(n389), .CPN(Clk_r), .Q(\Queue[4][0] ) );
  FDN1QM1P \Queue_reg[3][0]  ( .D(n517), .CPN(Clk_r), .Q(\Queue[3][0] ) );
  FDN1QM1P \Queue_reg[2][0]  ( .D(n485), .CPN(Clk_r), .Q(\Queue[2][0] ) );
  FDN1QM1P \Queue_reg[4][31]  ( .D(n388), .CPN(Clk_r), .Q(\Queue[4][31] ) );
  FDN1QM1P \Queue_reg[3][31]  ( .D(n548), .CPN(Clk_r), .Q(\Queue[3][31] ) );
  FDN1QM1P \Queue_reg[2][31]  ( .D(n516), .CPN(Clk_r), .Q(\Queue[2][31] ) );
  FDN2QM1P Full_reg ( .D(n420), .CPN(Clk_r), .CD(Rst_n), .Q(Full) );
  FDN1QM1P \Queue_reg[1][31]  ( .D(n452), .CPN(Clk_r), .Q(\Queue[1][31] ) );
  FDN1QM1P \Queue_reg[0][31]  ( .D(n484), .CPN(Clk_r), .Q(Packet_Out[31]) );
  FDN1QM1P \Queue_reg[1][30]  ( .D(n451), .CPN(Clk_r), .Q(\Queue[1][30] ) );
  FDN1QM1P \Queue_reg[0][30]  ( .D(n483), .CPN(Clk_r), .Q(Packet_Out[30]) );
  FDN1QM1P \Queue_reg[1][29]  ( .D(n450), .CPN(Clk_r), .Q(\Queue[1][29] ) );
  FDN1QM1P \Queue_reg[0][29]  ( .D(n482), .CPN(Clk_r), .Q(Packet_Out[29]) );
  FDN1QM1P \Queue_reg[1][28]  ( .D(n449), .CPN(Clk_r), .Q(\Queue[1][28] ) );
  FDN1QM1P \Queue_reg[0][28]  ( .D(n481), .CPN(Clk_r), .Q(Packet_Out[28]) );
  FDN1QM1P \Queue_reg[1][27]  ( .D(n448), .CPN(Clk_r), .Q(\Queue[1][27] ) );
  FDN1QM1P \Queue_reg[0][27]  ( .D(n480), .CPN(Clk_r), .Q(Packet_Out[27]) );
  FDN1QM1P \Queue_reg[1][26]  ( .D(n447), .CPN(Clk_r), .Q(\Queue[1][26] ) );
  FDN1QM1P \Queue_reg[0][26]  ( .D(n479), .CPN(Clk_r), .Q(Packet_Out[26]) );
  FDN1QM1P \Queue_reg[1][25]  ( .D(n446), .CPN(Clk_r), .Q(\Queue[1][25] ) );
  FDN1QM1P \Queue_reg[0][25]  ( .D(n478), .CPN(Clk_r), .Q(Packet_Out[25]) );
  FDN1QM1P \Queue_reg[1][24]  ( .D(n445), .CPN(Clk_r), .Q(\Queue[1][24] ) );
  FDN1QM1P \Queue_reg[0][24]  ( .D(n477), .CPN(Clk_r), .Q(Packet_Out[24]) );
  FDN1QM1P \Queue_reg[1][23]  ( .D(n444), .CPN(Clk_r), .Q(\Queue[1][23] ) );
  FDN1QM1P \Queue_reg[0][23]  ( .D(n476), .CPN(Clk_r), .Q(Packet_Out[23]) );
  FDN1QM1P \Queue_reg[1][22]  ( .D(n443), .CPN(Clk_r), .Q(\Queue[1][22] ) );
  FDN1QM1P \Queue_reg[0][22]  ( .D(n475), .CPN(Clk_r), .Q(Packet_Out[22]) );
  FDN1QM1P \Queue_reg[1][21]  ( .D(n442), .CPN(Clk_r), .Q(\Queue[1][21] ) );
  FDN1QM1P \Queue_reg[0][21]  ( .D(n474), .CPN(Clk_r), .Q(Packet_Out[21]) );
  FDN1QM1P \Queue_reg[1][20]  ( .D(n441), .CPN(Clk_r), .Q(\Queue[1][20] ) );
  FDN1QM1P \Queue_reg[0][20]  ( .D(n473), .CPN(Clk_r), .Q(Packet_Out[20]) );
  FDN1QM1P \Queue_reg[1][19]  ( .D(n440), .CPN(Clk_r), .Q(\Queue[1][19] ) );
  FDN1QM1P \Queue_reg[0][19]  ( .D(n472), .CPN(Clk_r), .Q(Packet_Out[19]) );
  FDN1QM1P \Queue_reg[1][18]  ( .D(n439), .CPN(Clk_r), .Q(\Queue[1][18] ) );
  FDN1QM1P \Queue_reg[0][18]  ( .D(n471), .CPN(Clk_r), .Q(Packet_Out[18]) );
  FDN1QM1P \Queue_reg[1][17]  ( .D(n438), .CPN(Clk_r), .Q(\Queue[1][17] ) );
  FDN1QM1P \Queue_reg[0][17]  ( .D(n470), .CPN(Clk_r), .Q(Packet_Out[17]) );
  FDN1QM1P \Queue_reg[1][16]  ( .D(n437), .CPN(Clk_r), .Q(\Queue[1][16] ) );
  FDN1QM1P \Queue_reg[0][16]  ( .D(n469), .CPN(Clk_r), .Q(Packet_Out[16]) );
  FDN1QM1P \Queue_reg[1][15]  ( .D(n436), .CPN(Clk_r), .Q(\Queue[1][15] ) );
  FDN1QM1P \Queue_reg[0][15]  ( .D(n468), .CPN(Clk_r), .Q(Packet_Out[15]) );
  FDN1QM1P \Queue_reg[1][14]  ( .D(n435), .CPN(Clk_r), .Q(\Queue[1][14] ) );
  FDN1QM1P \Queue_reg[0][14]  ( .D(n467), .CPN(Clk_r), .Q(Packet_Out[14]) );
  FDN1QM1P \Queue_reg[1][13]  ( .D(n434), .CPN(Clk_r), .Q(\Queue[1][13] ) );
  FDN1QM1P \Queue_reg[0][13]  ( .D(n466), .CPN(Clk_r), .Q(Packet_Out[13]) );
  FDN1QM1P \Queue_reg[1][12]  ( .D(n433), .CPN(Clk_r), .Q(\Queue[1][12] ) );
  FDN1QM1P \Queue_reg[0][12]  ( .D(n465), .CPN(Clk_r), .Q(Packet_Out[12]) );
  FDN1QM1P \Queue_reg[1][11]  ( .D(n432), .CPN(Clk_r), .Q(\Queue[1][11] ) );
  FDN1QM1P \Queue_reg[0][11]  ( .D(n464), .CPN(Clk_r), .Q(Packet_Out[11]) );
  FDN1QM1P \Queue_reg[1][10]  ( .D(n431), .CPN(Clk_r), .Q(\Queue[1][10] ) );
  FDN1QM1P \Queue_reg[0][10]  ( .D(n463), .CPN(Clk_r), .Q(Packet_Out[10]) );
  FDN1QM1P \Queue_reg[1][9]  ( .D(n430), .CPN(Clk_r), .Q(\Queue[1][9] ) );
  FDN1QM1P \Queue_reg[0][9]  ( .D(n462), .CPN(Clk_r), .Q(Packet_Out[9]) );
  FDN1QM1P \Queue_reg[1][8]  ( .D(n429), .CPN(Clk_r), .Q(\Queue[1][8] ) );
  FDN1QM1P \Queue_reg[0][8]  ( .D(n461), .CPN(Clk_r), .Q(Packet_Out[8]) );
  FDN1QM1P \Queue_reg[1][7]  ( .D(n428), .CPN(Clk_r), .Q(\Queue[1][7] ) );
  FDN1QM1P \Queue_reg[0][7]  ( .D(n460), .CPN(Clk_r), .Q(Packet_Out[7]) );
  FDN1QM1P \Queue_reg[1][6]  ( .D(n427), .CPN(Clk_r), .Q(\Queue[1][6] ) );
  FDN1QM1P \Queue_reg[0][6]  ( .D(n459), .CPN(Clk_r), .Q(Packet_Out[6]) );
  FDN1QM1P \Queue_reg[1][5]  ( .D(n426), .CPN(Clk_r), .Q(\Queue[1][5] ) );
  FDN1QM1P \Queue_reg[0][5]  ( .D(n458), .CPN(Clk_r), .Q(Packet_Out[5]) );
  FDN1QM1P \Queue_reg[1][4]  ( .D(n425), .CPN(Clk_r), .Q(\Queue[1][4] ) );
  FDN1QM1P \Queue_reg[0][4]  ( .D(n457), .CPN(Clk_r), .Q(Packet_Out[4]) );
  FDN1QM1P \Queue_reg[1][3]  ( .D(n424), .CPN(Clk_r), .Q(\Queue[1][3] ) );
  FDN1QM1P \Queue_reg[0][3]  ( .D(n456), .CPN(Clk_r), .Q(Packet_Out[3]) );
  FDN1QM1P \Queue_reg[1][2]  ( .D(n423), .CPN(Clk_r), .Q(\Queue[1][2] ) );
  FDN1QM1P \Queue_reg[0][2]  ( .D(n455), .CPN(Clk_r), .Q(Packet_Out[2]) );
  FDN1QM1P \Queue_reg[1][1]  ( .D(n422), .CPN(Clk_r), .Q(\Queue[1][1] ) );
  FDN1QM1P \Queue_reg[0][1]  ( .D(n454), .CPN(Clk_r), .Q(Packet_Out[1]) );
  FDN1QM1P \Queue_reg[1][0]  ( .D(n421), .CPN(Clk_r), .Q(\Queue[1][0] ) );
  FDN1QM1P \Queue_reg[0][0]  ( .D(n453), .CPN(Clk_r), .Q(Packet_Out[0]) );
  FDN2QM1P Empty_reg ( .D(n550), .CPN(Clk_r), .CD(Rst_n), .Q(n549) );
  BUFM2P U3 ( .A(n105), .Z(n11) );
  BUFM2P U4 ( .A(n140), .Z(n3) );
  N1M1P U5 ( .A(Read_Ack), .Z(n145) );
  ND2M1P U6 ( .A(Read_Ack), .B(Rst_n), .Z(n149) );
  N1M1P U7 ( .A(n4), .Z(n107) );
  OAI211M4P U8 ( .A(n108), .B(n145), .C(n4), .D(n32), .Z(n67) );
  NR2I1M8P U9 ( .A(n69), .B(n29), .Z(n28) );
  AOI21M3P U10 ( .A(n4), .B(n108), .C(n149), .Z(n65) );
  AOI21M3P U11 ( .A(n4), .B(n150), .C(n149), .Z(n377) );
  AOI21M3P U12 ( .A(n4), .B(n384), .C(n149), .Z(n103) );
  NR3M1P U13 ( .A(Count[2]), .B(n31), .C(n30), .Z(n148) );
  BUFM6P U14 ( .A(Write_Ack), .Z(n4) );
  BUFM2P U15 ( .A(n143), .Z(n16) );
  BUFM2P U16 ( .A(n380), .Z(n20) );
  BUFM2P U17 ( .A(n143), .Z(n15) );
  BUFM2P U18 ( .A(n380), .Z(n19) );
  OAI211M2P U19 ( .A(n148), .B(n145), .C(n4), .D(n106), .Z(n143) );
  OAI211M2P U20 ( .A(n150), .B(n145), .C(n4), .D(n144), .Z(n380) );
  OAI211M2P U21 ( .A(n148), .B(n147), .C(Rst_n), .D(n146), .Z(n378) );
  OAI211M2P U22 ( .A(n108), .B(n147), .C(Rst_n), .D(n146), .Z(n141) );
  ND2M1P U23 ( .A(n26), .B(Rst_n), .Z(n69) );
  N1M1P U24 ( .A(n150), .Z(n29) );
  NR2M2P U25 ( .A(Read_Ack), .B(n107), .Z(n26) );
  NR3M1P U26 ( .A(Count[0]), .B(Count[2]), .C(n30), .Z(n108) );
  NR3M1P U27 ( .A(Count[0]), .B(Count[1]), .C(n27), .Z(n150) );
  NR3M1P U28 ( .A(n31), .B(Count[2]), .C(Count[1]), .Z(n384) );
  N1M1P U29 ( .A(Count[0]), .Z(n31) );
  N1M1P U30 ( .A(Count[1]), .Z(n30) );
  N1M1P U31 ( .A(Count[2]), .Z(n27) );
  N1M1P U32 ( .A(Packet_In[23]), .Z(n198) );
  N1M1P U33 ( .A(Packet_In[25]), .Z(n202) );
  N1M1P U34 ( .A(Packet_In[29]), .Z(n374) );
  N1M1P U35 ( .A(Packet_In[27]), .Z(n206) );
  N1M1P U36 ( .A(Packet_In[28]), .Z(n208) );
  N1M1P U37 ( .A(Packet_In[26]), .Z(n204) );
  N1M1P U38 ( .A(Packet_In[31]), .Z(n381) );
  N1M1P U39 ( .A(Packet_In[24]), .Z(n200) );
  N1M1P U40 ( .A(Packet_In[22]), .Z(n196) );
  N1M1P U41 ( .A(Packet_In[21]), .Z(n194) );
  N1M1P U42 ( .A(Packet_In[20]), .Z(n192) );
  N1M1P U43 ( .A(Packet_In[9]), .Z(n170) );
  N1M1P U44 ( .A(Packet_In[30]), .Z(n376) );
  N1M1P U45 ( .A(Packet_In[13]), .Z(n178) );
  N1M1P U46 ( .A(Packet_In[7]), .Z(n166) );
  N1M1P U47 ( .A(Packet_In[14]), .Z(n180) );
  N1M1P U48 ( .A(Packet_In[17]), .Z(n186) );
  N1M1P U49 ( .A(Packet_In[12]), .Z(n176) );
  N1M1P U50 ( .A(Packet_In[19]), .Z(n190) );
  N1M1P U51 ( .A(Packet_In[11]), .Z(n174) );
  N1M1P U52 ( .A(Packet_In[18]), .Z(n188) );
  N1M1P U53 ( .A(Packet_In[15]), .Z(n182) );
  N1M1P U54 ( .A(Packet_In[16]), .Z(n184) );
  N1M1P U55 ( .A(Packet_In[10]), .Z(n172) );
  N1M1P U56 ( .A(Packet_In[8]), .Z(n168) );
  N1M1P U57 ( .A(Packet_In[1]), .Z(n154) );
  N1M1P U58 ( .A(Packet_In[6]), .Z(n164) );
  N1M1P U59 ( .A(Packet_In[5]), .Z(n162) );
  N1M1P U60 ( .A(Packet_In[4]), .Z(n160) );
  N1M1P U61 ( .A(Packet_In[3]), .Z(n158) );
  N1M1P U62 ( .A(Packet_In[2]), .Z(n156) );
  N1M1P U63 ( .A(Packet_In[0]), .Z(n152) );
  BUFM2P U64 ( .A(n105), .Z(n12) );
  BUFM2P U65 ( .A(n65), .Z(n8) );
  BUFM2P U66 ( .A(n141), .Z(n14) );
  BUFM2P U67 ( .A(n141), .Z(n13) );
  BUFM2P U68 ( .A(n378), .Z(n18) );
  BUFM2P U69 ( .A(n378), .Z(n17) );
  BUFM2P U70 ( .A(n64), .Z(n7) );
  BUFM2P U71 ( .A(n64), .Z(n6) );
  BUFM2P U72 ( .A(n64), .Z(n5) );
  N1M2P U73 ( .A(n26), .Z(n147) );
  BUFM2P U74 ( .A(n102), .Z(n10) );
  BUFM2P U75 ( .A(n102), .Z(n9) );
  N1M2P U76 ( .A(n70), .Z(n102) );
  OAI211M1P U77 ( .A(n384), .B(n145), .C(n4), .D(n70), .Z(n105) );
  NR2M1P U78 ( .A(n145), .B(n4), .Z(n383) );
  NR2M1P U79 ( .A(n26), .B(n383), .Z(n382) );
  AOI22CDNM1P U80 ( .A(n382), .B(n31), .C(n382), .D(n31), .Z(n385) );
  N1M1P U81 ( .A(n383), .Z(n25) );
  AOI22M1P U82 ( .A(Count[0]), .B(n147), .C(n25), .D(n31), .Z(n22) );
  AOI22CDNM1P U83 ( .A(Count[1]), .B(n22), .C(n22), .D(Count[1]), .Z(n386) );
  ND3M1P U84 ( .A(n31), .B(n27), .C(n30), .Z(n68) );
  ND2M1P U85 ( .A(Count[1]), .B(Read_Ack), .Z(n21) );
  OAI211M1P U86 ( .A(Count[1]), .B(n147), .C(n22), .D(n21), .Z(n23) );
  AOI22M1P U87 ( .A(n26), .B(n148), .C(Count[2]), .D(n23), .Z(n24) );
  OAI21M1P U88 ( .A(n68), .B(n25), .C(n24), .Z(n387) );
  AOI22CDNM1P U89 ( .A(n28), .B(n381), .C(\Queue[4][31] ), .D(n28), .Z(n388)
         );
  AOI22CDNM1P U90 ( .A(n28), .B(n152), .C(\Queue[4][0] ), .D(n28), .Z(n389) );
  AOI22CDNM1P U91 ( .A(n28), .B(n154), .C(\Queue[4][1] ), .D(n28), .Z(n390) );
  AOI22CDNM1P U92 ( .A(n28), .B(n156), .C(\Queue[4][2] ), .D(n28), .Z(n391) );
  AOI22CDNM1P U93 ( .A(n28), .B(n158), .C(\Queue[4][3] ), .D(n28), .Z(n392) );
  AOI22CDNM1P U94 ( .A(n28), .B(n160), .C(\Queue[4][4] ), .D(n28), .Z(n393) );
  AOI22CDNM1P U95 ( .A(n28), .B(n162), .C(\Queue[4][5] ), .D(n28), .Z(n394) );
  AOI22CDNM1P U96 ( .A(n28), .B(n164), .C(\Queue[4][6] ), .D(n28), .Z(n395) );
  AOI22CDNM1P U97 ( .A(n28), .B(n166), .C(\Queue[4][7] ), .D(n28), .Z(n396) );
  AOI22CDNM1P U98 ( .A(n28), .B(n168), .C(\Queue[4][8] ), .D(n28), .Z(n397) );
  AOI22CDNM1P U99 ( .A(n28), .B(n170), .C(\Queue[4][9] ), .D(n28), .Z(n398) );
  AOI22CDNM1P U100 ( .A(n28), .B(n172), .C(\Queue[4][10] ), .D(n28), .Z(n399)
         );
  AOI22CDNM1P U101 ( .A(n28), .B(n174), .C(\Queue[4][11] ), .D(n28), .Z(n400)
         );
  AOI22CDNM1P U102 ( .A(n28), .B(n176), .C(\Queue[4][12] ), .D(n28), .Z(n401)
         );
  AOI22CDNM1P U103 ( .A(n28), .B(n178), .C(\Queue[4][13] ), .D(n28), .Z(n402)
         );
  AOI22CDNM1P U104 ( .A(n28), .B(n180), .C(\Queue[4][14] ), .D(n28), .Z(n403)
         );
  AOI22CDNM1P U105 ( .A(n28), .B(n182), .C(\Queue[4][15] ), .D(n28), .Z(n404)
         );
  AOI22CDNM1P U106 ( .A(n28), .B(n184), .C(\Queue[4][16] ), .D(n28), .Z(n405)
         );
  AOI22CDNM1P U107 ( .A(n28), .B(n186), .C(\Queue[4][17] ), .D(n28), .Z(n406)
         );
  AOI22CDNM1P U108 ( .A(n28), .B(n188), .C(\Queue[4][18] ), .D(n28), .Z(n407)
         );
  AOI22CDNM1P U109 ( .A(n28), .B(n190), .C(\Queue[4][19] ), .D(n28), .Z(n408)
         );
  AOI22CDNM1P U110 ( .A(n28), .B(n192), .C(\Queue[4][20] ), .D(n28), .Z(n409)
         );
  AOI22CDNM1P U111 ( .A(n28), .B(n194), .C(\Queue[4][21] ), .D(n28), .Z(n410)
         );
  AOI22CDNM1P U112 ( .A(n28), .B(n196), .C(\Queue[4][22] ), .D(n28), .Z(n411)
         );
  AOI22CDNM1P U113 ( .A(n28), .B(n198), .C(\Queue[4][23] ), .D(n28), .Z(n412)
         );
  AOI22CDNM1P U114 ( .A(n28), .B(n200), .C(\Queue[4][24] ), .D(n28), .Z(n413)
         );
  AOI22CDNM1P U115 ( .A(n28), .B(n202), .C(\Queue[4][25] ), .D(n28), .Z(n414)
         );
  AOI22CDNM1P U116 ( .A(n28), .B(n204), .C(\Queue[4][26] ), .D(n28), .Z(n415)
         );
  AOI22CDNM1P U117 ( .A(n28), .B(n206), .C(\Queue[4][27] ), .D(n28), .Z(n416)
         );
  AOI22CDNM1P U118 ( .A(n28), .B(n208), .C(\Queue[4][28] ), .D(n28), .Z(n417)
         );
  AOI22CDNM1P U119 ( .A(n28), .B(n374), .C(\Queue[4][29] ), .D(n28), .Z(n418)
         );
  AOI22CDNM1P U120 ( .A(n28), .B(n376), .C(\Queue[4][30] ), .D(n28), .Z(n419)
         );
  OAI22CDNM1P U121 ( .A(n147), .B(n29), .C(n382), .D(Full), .Z(n420) );
  OA21M1P U122 ( .A(n147), .B(n384), .C(Rst_n), .Z(n32) );
  OAI21M1P U123 ( .A(n4), .B(Read_Ack), .C(n32), .Z(n64) );
  AOI22M1P U124 ( .A(\Queue[2][0] ), .B(n65), .C(\Queue[1][0] ), .D(n5), .Z(
        n33) );
  OAI21M1P U125 ( .A(n152), .B(n67), .C(n33), .Z(n421) );
  AOI22M1P U126 ( .A(n8), .B(\Queue[2][1] ), .C(\Queue[1][1] ), .D(n5), .Z(n34) );
  OAI21M1P U127 ( .A(n67), .B(n154), .C(n34), .Z(n422) );
  AOI22M1P U128 ( .A(n65), .B(\Queue[2][2] ), .C(\Queue[1][2] ), .D(n5), .Z(
        n35) );
  OAI21M1P U129 ( .A(n67), .B(n156), .C(n35), .Z(n423) );
  AOI22M1P U130 ( .A(n65), .B(\Queue[2][3] ), .C(\Queue[1][3] ), .D(n5), .Z(
        n36) );
  OAI21M1P U131 ( .A(n67), .B(n158), .C(n36), .Z(n424) );
  AOI22M1P U132 ( .A(n65), .B(\Queue[2][4] ), .C(\Queue[1][4] ), .D(n5), .Z(
        n37) );
  OAI21M1P U133 ( .A(n67), .B(n160), .C(n37), .Z(n425) );
  AOI22M1P U134 ( .A(n65), .B(\Queue[2][5] ), .C(\Queue[1][5] ), .D(n5), .Z(
        n38) );
  OAI21M1P U135 ( .A(n67), .B(n162), .C(n38), .Z(n426) );
  AOI22M1P U136 ( .A(n65), .B(\Queue[2][6] ), .C(\Queue[1][6] ), .D(n5), .Z(
        n39) );
  OAI21M1P U137 ( .A(n67), .B(n164), .C(n39), .Z(n427) );
  AOI22M1P U138 ( .A(n65), .B(\Queue[2][7] ), .C(\Queue[1][7] ), .D(n5), .Z(
        n40) );
  OAI21M1P U139 ( .A(n67), .B(n166), .C(n40), .Z(n428) );
  AOI22M1P U140 ( .A(n65), .B(\Queue[2][8] ), .C(\Queue[1][8] ), .D(n5), .Z(
        n41) );
  OAI21M1P U141 ( .A(n67), .B(n168), .C(n41), .Z(n429) );
  AOI22M1P U142 ( .A(n65), .B(\Queue[2][9] ), .C(\Queue[1][9] ), .D(n6), .Z(
        n42) );
  OAI21M1P U143 ( .A(n67), .B(n170), .C(n42), .Z(n430) );
  AOI22M1P U144 ( .A(n65), .B(\Queue[2][10] ), .C(\Queue[1][10] ), .D(n6), .Z(
        n43) );
  OAI21M1P U145 ( .A(n67), .B(n172), .C(n43), .Z(n431) );
  AOI22M1P U146 ( .A(n65), .B(\Queue[2][11] ), .C(\Queue[1][11] ), .D(n6), .Z(
        n44) );
  OAI21M1P U147 ( .A(n67), .B(n174), .C(n44), .Z(n432) );
  AOI22M1P U148 ( .A(n8), .B(\Queue[2][12] ), .C(\Queue[1][12] ), .D(n6), .Z(
        n45) );
  OAI21M1P U149 ( .A(n67), .B(n176), .C(n45), .Z(n433) );
  AOI22M1P U150 ( .A(n8), .B(\Queue[2][13] ), .C(\Queue[1][13] ), .D(n6), .Z(
        n46) );
  OAI21M1P U151 ( .A(n67), .B(n178), .C(n46), .Z(n434) );
  AOI22M1P U152 ( .A(n8), .B(\Queue[2][14] ), .C(\Queue[1][14] ), .D(n6), .Z(
        n47) );
  OAI21M1P U153 ( .A(n67), .B(n180), .C(n47), .Z(n435) );
  AOI22M1P U154 ( .A(n8), .B(\Queue[2][15] ), .C(\Queue[1][15] ), .D(n6), .Z(
        n48) );
  OAI21M1P U155 ( .A(n67), .B(n182), .C(n48), .Z(n436) );
  AOI22M1P U156 ( .A(n8), .B(\Queue[2][16] ), .C(\Queue[1][16] ), .D(n6), .Z(
        n49) );
  OAI21M1P U157 ( .A(n67), .B(n184), .C(n49), .Z(n437) );
  AOI22M1P U158 ( .A(n8), .B(\Queue[2][17] ), .C(\Queue[1][17] ), .D(n6), .Z(
        n50) );
  OAI21M1P U159 ( .A(n67), .B(n186), .C(n50), .Z(n438) );
  AOI22M1P U160 ( .A(n8), .B(\Queue[2][18] ), .C(\Queue[1][18] ), .D(n7), .Z(
        n51) );
  OAI21M1P U161 ( .A(n67), .B(n188), .C(n51), .Z(n439) );
  AOI22M1P U162 ( .A(n8), .B(\Queue[2][19] ), .C(\Queue[1][19] ), .D(n7), .Z(
        n52) );
  OAI21M1P U163 ( .A(n67), .B(n190), .C(n52), .Z(n440) );
  AOI22M1P U164 ( .A(n8), .B(\Queue[2][20] ), .C(\Queue[1][20] ), .D(n7), .Z(
        n53) );
  OAI21M1P U165 ( .A(n67), .B(n192), .C(n53), .Z(n441) );
  AOI22M1P U166 ( .A(n8), .B(\Queue[2][21] ), .C(\Queue[1][21] ), .D(n7), .Z(
        n54) );
  OAI21M1P U167 ( .A(n67), .B(n194), .C(n54), .Z(n442) );
  AOI22M1P U168 ( .A(n8), .B(\Queue[2][22] ), .C(\Queue[1][22] ), .D(n7), .Z(
        n55) );
  OAI21M1P U169 ( .A(n67), .B(n196), .C(n55), .Z(n443) );
  AOI22M1P U170 ( .A(n8), .B(\Queue[2][23] ), .C(\Queue[1][23] ), .D(n7), .Z(
        n56) );
  OAI21M1P U171 ( .A(n67), .B(n198), .C(n56), .Z(n444) );
  AOI22M1P U172 ( .A(n65), .B(\Queue[2][24] ), .C(\Queue[1][24] ), .D(n7), .Z(
        n57) );
  OAI21M1P U173 ( .A(n67), .B(n200), .C(n57), .Z(n445) );
  AOI22M1P U174 ( .A(n65), .B(\Queue[2][25] ), .C(\Queue[1][25] ), .D(n7), .Z(
        n58) );
  OAI21M1P U175 ( .A(n67), .B(n202), .C(n58), .Z(n446) );
  AOI22M1P U176 ( .A(n65), .B(\Queue[2][26] ), .C(\Queue[1][26] ), .D(n7), .Z(
        n59) );
  OAI21M1P U177 ( .A(n67), .B(n204), .C(n59), .Z(n447) );
  AOI22M1P U178 ( .A(n65), .B(\Queue[2][27] ), .C(\Queue[1][27] ), .D(n7), .Z(
        n60) );
  OAI21M1P U179 ( .A(n67), .B(n206), .C(n60), .Z(n448) );
  AOI22M1P U180 ( .A(n65), .B(\Queue[2][28] ), .C(\Queue[1][28] ), .D(n5), .Z(
        n61) );
  OAI21M1P U181 ( .A(n67), .B(n208), .C(n61), .Z(n449) );
  AOI22M1P U182 ( .A(n65), .B(\Queue[2][29] ), .C(\Queue[1][29] ), .D(n6), .Z(
        n62) );
  OAI21M1P U183 ( .A(n67), .B(n374), .C(n62), .Z(n450) );
  AOI22M1P U184 ( .A(n65), .B(\Queue[2][30] ), .C(\Queue[1][30] ), .D(n7), .Z(
        n63) );
  OAI21M1P U185 ( .A(n67), .B(n376), .C(n63), .Z(n451) );
  AOI22M1P U186 ( .A(n65), .B(\Queue[2][31] ), .C(\Queue[1][31] ), .D(n5), .Z(
        n66) );
  OAI21M1P U187 ( .A(n67), .B(n381), .C(n66), .Z(n452) );
  OAI21M1P U188 ( .A(n69), .B(n68), .C(n149), .Z(n70) );
  AOI22M1P U189 ( .A(\Queue[1][0] ), .B(n103), .C(n9), .D(Packet_Out[0]), .Z(
        n71) );
  OAI21M1P U190 ( .A(n152), .B(n11), .C(n71), .Z(n453) );
  AOI22M1P U191 ( .A(\Queue[1][1] ), .B(n103), .C(n9), .D(Packet_Out[1]), .Z(
        n72) );
  OAI21M1P U192 ( .A(n154), .B(n11), .C(n72), .Z(n454) );
  AOI22M1P U193 ( .A(\Queue[1][2] ), .B(n103), .C(n9), .D(Packet_Out[2]), .Z(
        n73) );
  OAI21M1P U194 ( .A(n156), .B(n11), .C(n73), .Z(n455) );
  AOI22M1P U195 ( .A(\Queue[1][3] ), .B(n103), .C(n9), .D(Packet_Out[3]), .Z(
        n74) );
  OAI21M1P U196 ( .A(n158), .B(n11), .C(n74), .Z(n456) );
  AOI22M1P U197 ( .A(\Queue[1][4] ), .B(n103), .C(n9), .D(Packet_Out[4]), .Z(
        n75) );
  OAI21M1P U198 ( .A(n160), .B(n11), .C(n75), .Z(n457) );
  AOI22M1P U199 ( .A(\Queue[1][5] ), .B(n103), .C(n9), .D(Packet_Out[5]), .Z(
        n76) );
  OAI21M1P U200 ( .A(n162), .B(n11), .C(n76), .Z(n458) );
  AOI22M1P U201 ( .A(\Queue[1][6] ), .B(n103), .C(n9), .D(Packet_Out[6]), .Z(
        n77) );
  OAI21M1P U202 ( .A(n164), .B(n11), .C(n77), .Z(n459) );
  AOI22M1P U203 ( .A(\Queue[1][7] ), .B(n103), .C(n9), .D(Packet_Out[7]), .Z(
        n78) );
  OAI21M1P U204 ( .A(n166), .B(n11), .C(n78), .Z(n460) );
  AOI22M1P U205 ( .A(\Queue[1][8] ), .B(n103), .C(n9), .D(Packet_Out[8]), .Z(
        n79) );
  OAI21M1P U206 ( .A(n168), .B(n11), .C(n79), .Z(n461) );
  AOI22M1P U207 ( .A(\Queue[1][9] ), .B(n103), .C(n9), .D(Packet_Out[9]), .Z(
        n80) );
  OAI21M1P U208 ( .A(n170), .B(n11), .C(n80), .Z(n462) );
  AOI22M1P U209 ( .A(\Queue[1][10] ), .B(n103), .C(n102), .D(Packet_Out[10]), 
        .Z(n81) );
  OAI21M1P U210 ( .A(n172), .B(n11), .C(n81), .Z(n463) );
  AOI22M1P U211 ( .A(\Queue[1][11] ), .B(n103), .C(n102), .D(Packet_Out[11]), 
        .Z(n82) );
  OAI21M1P U212 ( .A(n174), .B(n11), .C(n82), .Z(n464) );
  AOI22M1P U213 ( .A(\Queue[1][12] ), .B(n103), .C(n102), .D(Packet_Out[12]), 
        .Z(n83) );
  OAI21M1P U214 ( .A(n176), .B(n11), .C(n83), .Z(n465) );
  AOI22M1P U215 ( .A(\Queue[1][13] ), .B(n103), .C(n102), .D(Packet_Out[13]), 
        .Z(n84) );
  OAI21M1P U216 ( .A(n178), .B(n11), .C(n84), .Z(n466) );
  AOI22M1P U217 ( .A(\Queue[1][14] ), .B(n103), .C(n102), .D(Packet_Out[14]), 
        .Z(n85) );
  OAI21M1P U218 ( .A(n180), .B(n11), .C(n85), .Z(n467) );
  AOI22M1P U219 ( .A(\Queue[1][15] ), .B(n103), .C(n102), .D(Packet_Out[15]), 
        .Z(n86) );
  OAI21M1P U220 ( .A(n182), .B(n11), .C(n86), .Z(n468) );
  AOI22M1P U221 ( .A(\Queue[1][16] ), .B(n103), .C(n102), .D(Packet_Out[16]), 
        .Z(n87) );
  OAI21M1P U222 ( .A(n184), .B(n11), .C(n87), .Z(n469) );
  AOI22M1P U223 ( .A(\Queue[1][17] ), .B(n103), .C(n102), .D(Packet_Out[17]), 
        .Z(n88) );
  OAI21M1P U224 ( .A(n186), .B(n11), .C(n88), .Z(n470) );
  AOI22M1P U225 ( .A(\Queue[1][18] ), .B(n103), .C(n102), .D(Packet_Out[18]), 
        .Z(n89) );
  OAI21M1P U226 ( .A(n188), .B(n11), .C(n89), .Z(n471) );
  AOI22M1P U227 ( .A(\Queue[1][19] ), .B(n103), .C(n102), .D(Packet_Out[19]), 
        .Z(n90) );
  OAI21M1P U228 ( .A(n190), .B(n11), .C(n90), .Z(n472) );
  AOI22M1P U229 ( .A(\Queue[1][20] ), .B(n103), .C(n10), .D(Packet_Out[20]), 
        .Z(n91) );
  OAI21M1P U230 ( .A(n192), .B(n12), .C(n91), .Z(n473) );
  AOI22M1P U231 ( .A(\Queue[1][21] ), .B(n103), .C(n10), .D(Packet_Out[21]), 
        .Z(n92) );
  OAI21M1P U232 ( .A(n194), .B(n12), .C(n92), .Z(n474) );
  AOI22M1P U233 ( .A(\Queue[1][22] ), .B(n103), .C(n10), .D(Packet_Out[22]), 
        .Z(n93) );
  OAI21M1P U234 ( .A(n196), .B(n12), .C(n93), .Z(n475) );
  AOI22M1P U235 ( .A(\Queue[1][23] ), .B(n103), .C(n10), .D(Packet_Out[23]), 
        .Z(n94) );
  OAI21M1P U236 ( .A(n198), .B(n12), .C(n94), .Z(n476) );
  AOI22M1P U237 ( .A(\Queue[1][24] ), .B(n103), .C(n10), .D(Packet_Out[24]), 
        .Z(n95) );
  OAI21M1P U238 ( .A(n200), .B(n12), .C(n95), .Z(n477) );
  AOI22M1P U239 ( .A(\Queue[1][25] ), .B(n103), .C(n10), .D(Packet_Out[25]), 
        .Z(n96) );
  OAI21M1P U240 ( .A(n202), .B(n12), .C(n96), .Z(n478) );
  AOI22M1P U241 ( .A(\Queue[1][26] ), .B(n103), .C(n10), .D(Packet_Out[26]), 
        .Z(n97) );
  OAI21M1P U242 ( .A(n204), .B(n12), .C(n97), .Z(n479) );
  AOI22M1P U243 ( .A(\Queue[1][27] ), .B(n103), .C(n10), .D(Packet_Out[27]), 
        .Z(n98) );
  OAI21M1P U244 ( .A(n206), .B(n12), .C(n98), .Z(n480) );
  AOI22M1P U245 ( .A(\Queue[1][28] ), .B(n103), .C(n10), .D(Packet_Out[28]), 
        .Z(n99) );
  OAI21M1P U246 ( .A(n208), .B(n12), .C(n99), .Z(n481) );
  AOI22M1P U247 ( .A(\Queue[1][29] ), .B(n103), .C(n10), .D(Packet_Out[29]), 
        .Z(n100) );
  OAI21M1P U248 ( .A(n374), .B(n12), .C(n100), .Z(n482) );
  AOI22M1P U249 ( .A(\Queue[1][30] ), .B(n103), .C(n10), .D(Packet_Out[30]), 
        .Z(n101) );
  OAI21M1P U250 ( .A(n376), .B(n11), .C(n101), .Z(n483) );
  AOI22M1P U251 ( .A(\Queue[1][31] ), .B(n103), .C(n9), .D(Packet_Out[31]), 
        .Z(n104) );
  OAI21M1P U252 ( .A(n381), .B(n12), .C(n104), .Z(n484) );
  OA21M1P U253 ( .A(n147), .B(n108), .C(Rst_n), .Z(n106) );
  ND2M1P U254 ( .A(n107), .B(n145), .Z(n146) );
  AOI21M1P U255 ( .A(n4), .B(n148), .C(n149), .Z(n140) );
  AOI22M1P U256 ( .A(\Queue[2][0] ), .B(n141), .C(\Queue[3][0] ), .D(n3), .Z(
        n109) );
  OAI21M1P U257 ( .A(n152), .B(n16), .C(n109), .Z(n485) );
  AOI22M1P U258 ( .A(\Queue[2][1] ), .B(n141), .C(n3), .D(\Queue[3][1] ), .Z(
        n110) );
  OAI21M1P U259 ( .A(n154), .B(n143), .C(n110), .Z(n486) );
  AOI22M1P U260 ( .A(\Queue[2][2] ), .B(n141), .C(n3), .D(\Queue[3][2] ), .Z(
        n111) );
  OAI21M1P U261 ( .A(n156), .B(n143), .C(n111), .Z(n487) );
  AOI22M1P U262 ( .A(\Queue[2][3] ), .B(n141), .C(n3), .D(\Queue[3][3] ), .Z(
        n112) );
  OAI21M1P U263 ( .A(n158), .B(n143), .C(n112), .Z(n488) );
  AOI22M1P U264 ( .A(\Queue[2][4] ), .B(n141), .C(n3), .D(\Queue[3][4] ), .Z(
        n113) );
  OAI21M1P U265 ( .A(n160), .B(n143), .C(n113), .Z(n489) );
  AOI22M1P U266 ( .A(\Queue[2][5] ), .B(n141), .C(n3), .D(\Queue[3][5] ), .Z(
        n114) );
  OAI21M1P U267 ( .A(n162), .B(n143), .C(n114), .Z(n490) );
  AOI22M1P U268 ( .A(\Queue[2][6] ), .B(n13), .C(n3), .D(\Queue[3][6] ), .Z(
        n115) );
  OAI21M1P U269 ( .A(n164), .B(n143), .C(n115), .Z(n491) );
  AOI22M1P U270 ( .A(\Queue[2][7] ), .B(n14), .C(n3), .D(\Queue[3][7] ), .Z(
        n116) );
  OAI21M1P U271 ( .A(n166), .B(n15), .C(n116), .Z(n492) );
  AOI22M1P U272 ( .A(\Queue[2][8] ), .B(n13), .C(n3), .D(\Queue[3][8] ), .Z(
        n117) );
  OAI21M1P U273 ( .A(n168), .B(n16), .C(n117), .Z(n493) );
  AOI22M1P U274 ( .A(\Queue[2][9] ), .B(n14), .C(n3), .D(\Queue[3][9] ), .Z(
        n118) );
  OAI21M1P U275 ( .A(n170), .B(n15), .C(n118), .Z(n494) );
  AOI22M1P U276 ( .A(\Queue[2][10] ), .B(n13), .C(n3), .D(\Queue[3][10] ), .Z(
        n119) );
  OAI21M1P U277 ( .A(n172), .B(n15), .C(n119), .Z(n495) );
  AOI22M1P U278 ( .A(\Queue[2][11] ), .B(n13), .C(n3), .D(\Queue[3][11] ), .Z(
        n120) );
  OAI21M1P U279 ( .A(n174), .B(n15), .C(n120), .Z(n496) );
  AOI22M1P U280 ( .A(\Queue[2][12] ), .B(n13), .C(n3), .D(\Queue[3][12] ), .Z(
        n121) );
  OAI21M1P U281 ( .A(n176), .B(n15), .C(n121), .Z(n497) );
  AOI22M1P U282 ( .A(\Queue[2][13] ), .B(n13), .C(n3), .D(\Queue[3][13] ), .Z(
        n122) );
  OAI21M1P U283 ( .A(n178), .B(n15), .C(n122), .Z(n498) );
  AOI22M1P U284 ( .A(\Queue[2][14] ), .B(n13), .C(n3), .D(\Queue[3][14] ), .Z(
        n123) );
  OAI21M1P U285 ( .A(n180), .B(n15), .C(n123), .Z(n499) );
  AOI22M1P U286 ( .A(\Queue[2][15] ), .B(n13), .C(n3), .D(\Queue[3][15] ), .Z(
        n124) );
  OAI21M1P U287 ( .A(n182), .B(n15), .C(n124), .Z(n500) );
  AOI22M1P U288 ( .A(\Queue[2][16] ), .B(n13), .C(n3), .D(\Queue[3][16] ), .Z(
        n125) );
  OAI21M1P U289 ( .A(n184), .B(n15), .C(n125), .Z(n501) );
  AOI22M1P U290 ( .A(\Queue[2][17] ), .B(n13), .C(n3), .D(\Queue[3][17] ), .Z(
        n126) );
  OAI21M1P U291 ( .A(n186), .B(n15), .C(n126), .Z(n502) );
  AOI22M1P U292 ( .A(\Queue[2][18] ), .B(n13), .C(n3), .D(\Queue[3][18] ), .Z(
        n127) );
  OAI21M1P U293 ( .A(n188), .B(n15), .C(n127), .Z(n503) );
  AOI22M1P U294 ( .A(\Queue[2][19] ), .B(n13), .C(n3), .D(\Queue[3][19] ), .Z(
        n128) );
  OAI21M1P U295 ( .A(n190), .B(n15), .C(n128), .Z(n504) );
  AOI22M1P U296 ( .A(\Queue[2][20] ), .B(n14), .C(n3), .D(\Queue[3][20] ), .Z(
        n129) );
  OAI21M1P U297 ( .A(n192), .B(n16), .C(n129), .Z(n505) );
  AOI22M1P U298 ( .A(\Queue[2][21] ), .B(n14), .C(n3), .D(\Queue[3][21] ), .Z(
        n130) );
  OAI21M1P U299 ( .A(n194), .B(n16), .C(n130), .Z(n506) );
  AOI22M1P U300 ( .A(\Queue[2][22] ), .B(n14), .C(n3), .D(\Queue[3][22] ), .Z(
        n131) );
  OAI21M1P U301 ( .A(n196), .B(n16), .C(n131), .Z(n507) );
  AOI22M1P U302 ( .A(\Queue[2][23] ), .B(n14), .C(n3), .D(\Queue[3][23] ), .Z(
        n132) );
  OAI21M1P U303 ( .A(n198), .B(n16), .C(n132), .Z(n508) );
  AOI22M1P U304 ( .A(\Queue[2][24] ), .B(n14), .C(n3), .D(\Queue[3][24] ), .Z(
        n133) );
  OAI21M1P U305 ( .A(n200), .B(n16), .C(n133), .Z(n509) );
  AOI22M1P U306 ( .A(\Queue[2][25] ), .B(n14), .C(n3), .D(\Queue[3][25] ), .Z(
        n134) );
  OAI21M1P U307 ( .A(n202), .B(n16), .C(n134), .Z(n510) );
  AOI22M1P U308 ( .A(\Queue[2][26] ), .B(n14), .C(n3), .D(\Queue[3][26] ), .Z(
        n135) );
  OAI21M1P U309 ( .A(n204), .B(n16), .C(n135), .Z(n511) );
  AOI22M1P U310 ( .A(\Queue[2][27] ), .B(n14), .C(n3), .D(\Queue[3][27] ), .Z(
        n136) );
  OAI21M1P U311 ( .A(n206), .B(n16), .C(n136), .Z(n512) );
  AOI22M1P U312 ( .A(\Queue[2][28] ), .B(n14), .C(n3), .D(\Queue[3][28] ), .Z(
        n137) );
  OAI21M1P U313 ( .A(n208), .B(n16), .C(n137), .Z(n513) );
  AOI22M1P U314 ( .A(\Queue[2][29] ), .B(n14), .C(n3), .D(\Queue[3][29] ), .Z(
        n138) );
  OAI21M1P U315 ( .A(n374), .B(n16), .C(n138), .Z(n514) );
  AOI22M1P U316 ( .A(\Queue[2][30] ), .B(n13), .C(n3), .D(\Queue[3][30] ), .Z(
        n139) );
  OAI21M1P U317 ( .A(n376), .B(n15), .C(n139), .Z(n515) );
  AOI22M1P U318 ( .A(\Queue[2][31] ), .B(n14), .C(n3), .D(\Queue[3][31] ), .Z(
        n142) );
  OAI21M1P U319 ( .A(n381), .B(n16), .C(n142), .Z(n516) );
  OA21M1P U320 ( .A(n147), .B(n148), .C(Rst_n), .Z(n144) );
  AOI22M1P U321 ( .A(\Queue[3][0] ), .B(n18), .C(n377), .D(\Queue[4][0] ), .Z(
        n151) );
  OAI21M1P U322 ( .A(n152), .B(n20), .C(n151), .Z(n517) );
  AOI22M1P U323 ( .A(\Queue[3][1] ), .B(n378), .C(n377), .D(\Queue[4][1] ), 
        .Z(n153) );
  OAI21M1P U324 ( .A(n154), .B(n380), .C(n153), .Z(n518) );
  AOI22M1P U325 ( .A(\Queue[3][2] ), .B(n378), .C(n377), .D(\Queue[4][2] ), 
        .Z(n155) );
  OAI21M1P U326 ( .A(n156), .B(n380), .C(n155), .Z(n519) );
  AOI22M1P U327 ( .A(\Queue[3][3] ), .B(n378), .C(n377), .D(\Queue[4][3] ), 
        .Z(n157) );
  OAI21M1P U328 ( .A(n158), .B(n380), .C(n157), .Z(n520) );
  AOI22M1P U329 ( .A(\Queue[3][4] ), .B(n378), .C(n377), .D(\Queue[4][4] ), 
        .Z(n159) );
  OAI21M1P U330 ( .A(n160), .B(n380), .C(n159), .Z(n521) );
  AOI22M1P U331 ( .A(\Queue[3][5] ), .B(n378), .C(n377), .D(\Queue[4][5] ), 
        .Z(n161) );
  OAI21M1P U332 ( .A(n162), .B(n380), .C(n161), .Z(n522) );
  AOI22M1P U333 ( .A(\Queue[3][6] ), .B(n378), .C(n377), .D(\Queue[4][6] ), 
        .Z(n163) );
  OAI21M1P U334 ( .A(n164), .B(n380), .C(n163), .Z(n523) );
  AOI22M1P U335 ( .A(\Queue[3][7] ), .B(n17), .C(n377), .D(\Queue[4][7] ), .Z(
        n165) );
  OAI21M1P U336 ( .A(n166), .B(n19), .C(n165), .Z(n524) );
  AOI22M1P U337 ( .A(\Queue[3][8] ), .B(n18), .C(n377), .D(\Queue[4][8] ), .Z(
        n167) );
  OAI21M1P U338 ( .A(n168), .B(n20), .C(n167), .Z(n525) );
  AOI22M1P U339 ( .A(\Queue[3][9] ), .B(n17), .C(n377), .D(\Queue[4][9] ), .Z(
        n169) );
  OAI21M1P U340 ( .A(n170), .B(n19), .C(n169), .Z(n526) );
  AOI22M1P U341 ( .A(\Queue[3][10] ), .B(n17), .C(n377), .D(\Queue[4][10] ), 
        .Z(n171) );
  OAI21M1P U342 ( .A(n172), .B(n19), .C(n171), .Z(n527) );
  AOI22M1P U343 ( .A(\Queue[3][11] ), .B(n17), .C(n377), .D(\Queue[4][11] ), 
        .Z(n173) );
  OAI21M1P U344 ( .A(n174), .B(n19), .C(n173), .Z(n528) );
  AOI22M1P U345 ( .A(\Queue[3][12] ), .B(n17), .C(n377), .D(\Queue[4][12] ), 
        .Z(n175) );
  OAI21M1P U346 ( .A(n176), .B(n19), .C(n175), .Z(n529) );
  AOI22M1P U347 ( .A(\Queue[3][13] ), .B(n17), .C(n377), .D(\Queue[4][13] ), 
        .Z(n177) );
  OAI21M1P U348 ( .A(n178), .B(n19), .C(n177), .Z(n530) );
  AOI22M1P U349 ( .A(\Queue[3][14] ), .B(n17), .C(n377), .D(\Queue[4][14] ), 
        .Z(n179) );
  OAI21M1P U350 ( .A(n180), .B(n19), .C(n179), .Z(n531) );
  AOI22M1P U351 ( .A(\Queue[3][15] ), .B(n17), .C(n377), .D(\Queue[4][15] ), 
        .Z(n181) );
  OAI21M1P U352 ( .A(n182), .B(n19), .C(n181), .Z(n532) );
  AOI22M1P U353 ( .A(\Queue[3][16] ), .B(n17), .C(n377), .D(\Queue[4][16] ), 
        .Z(n183) );
  OAI21M1P U354 ( .A(n184), .B(n19), .C(n183), .Z(n533) );
  AOI22M1P U355 ( .A(\Queue[3][17] ), .B(n17), .C(n377), .D(\Queue[4][17] ), 
        .Z(n185) );
  OAI21M1P U356 ( .A(n186), .B(n19), .C(n185), .Z(n534) );
  AOI22M1P U357 ( .A(\Queue[3][18] ), .B(n17), .C(n377), .D(\Queue[4][18] ), 
        .Z(n187) );
  OAI21M1P U358 ( .A(n188), .B(n19), .C(n187), .Z(n535) );
  AOI22M1P U359 ( .A(\Queue[3][19] ), .B(n17), .C(n377), .D(\Queue[4][19] ), 
        .Z(n189) );
  OAI21M1P U360 ( .A(n190), .B(n19), .C(n189), .Z(n536) );
  AOI22M1P U361 ( .A(\Queue[3][20] ), .B(n18), .C(n377), .D(\Queue[4][20] ), 
        .Z(n191) );
  OAI21M1P U362 ( .A(n192), .B(n20), .C(n191), .Z(n537) );
  AOI22M1P U363 ( .A(\Queue[3][21] ), .B(n18), .C(n377), .D(\Queue[4][21] ), 
        .Z(n193) );
  OAI21M1P U364 ( .A(n194), .B(n20), .C(n193), .Z(n538) );
  AOI22M1P U365 ( .A(\Queue[3][22] ), .B(n18), .C(n377), .D(\Queue[4][22] ), 
        .Z(n195) );
  OAI21M1P U366 ( .A(n196), .B(n20), .C(n195), .Z(n539) );
  AOI22M1P U367 ( .A(\Queue[3][23] ), .B(n18), .C(n377), .D(\Queue[4][23] ), 
        .Z(n197) );
  OAI21M1P U368 ( .A(n198), .B(n20), .C(n197), .Z(n540) );
  AOI22M1P U369 ( .A(\Queue[3][24] ), .B(n18), .C(n377), .D(\Queue[4][24] ), 
        .Z(n199) );
  OAI21M1P U370 ( .A(n200), .B(n20), .C(n199), .Z(n541) );
  AOI22M1P U371 ( .A(\Queue[3][25] ), .B(n18), .C(n377), .D(\Queue[4][25] ), 
        .Z(n201) );
  OAI21M1P U372 ( .A(n202), .B(n20), .C(n201), .Z(n542) );
  AOI22M1P U373 ( .A(\Queue[3][26] ), .B(n18), .C(n377), .D(\Queue[4][26] ), 
        .Z(n203) );
  OAI21M1P U374 ( .A(n204), .B(n20), .C(n203), .Z(n543) );
  AOI22M1P U375 ( .A(\Queue[3][27] ), .B(n18), .C(n377), .D(\Queue[4][27] ), 
        .Z(n205) );
  OAI21M1P U376 ( .A(n206), .B(n20), .C(n205), .Z(n544) );
  AOI22M1P U377 ( .A(\Queue[3][28] ), .B(n18), .C(n377), .D(\Queue[4][28] ), 
        .Z(n207) );
  OAI21M1P U378 ( .A(n208), .B(n20), .C(n207), .Z(n545) );
  AOI22M1P U379 ( .A(\Queue[3][29] ), .B(n18), .C(n377), .D(\Queue[4][29] ), 
        .Z(n373) );
  OAI21M1P U380 ( .A(n374), .B(n20), .C(n373), .Z(n546) );
  AOI22M1P U381 ( .A(\Queue[3][30] ), .B(n17), .C(n377), .D(\Queue[4][30] ), 
        .Z(n375) );
  OAI21M1P U382 ( .A(n376), .B(n19), .C(n375), .Z(n547) );
  AOI22M1P U383 ( .A(\Queue[3][31] ), .B(n18), .C(n377), .D(\Queue[4][31] ), 
        .Z(n379) );
  OAI21M1P U384 ( .A(n381), .B(n20), .C(n379), .Z(n548) );
  N1M1P U385 ( .A(n549), .Z(Empty) );
  AOI22M1P U386 ( .A(n384), .B(n383), .C(n382), .D(Empty), .Z(n550) );
endmodule


module Link_Control_1 ( Clk_r, Rst_n, Tx_Ready, Tx_Error, RxData_Valid, RxData, 
        Packet_From_Core, TxQueue_Write, RxQueue_Read, TxData_Valid, TxData, 
        Error_Ack, Core_Rcv_Ready, Packet_To_Core, RxQueue_Empty, TxQueue_Full
 );
  input [31:0] RxData;
  input [31:0] Packet_From_Core;
  output [31:0] TxData;
  output [31:0] Packet_To_Core;
  input Clk_r, Rst_n, Tx_Ready, Tx_Error, RxData_Valid, TxQueue_Write,
         RxQueue_Read;
  output TxData_Valid, Error_Ack, Core_Rcv_Ready, RxQueue_Empty, TxQueue_Full;
  wire   TxQueue_Read, TxQueue_Empty, RxQueue_Write, RxQueue_Full, N9, N16, n5,
         n6, n7, n8, n9;

  Packet_Queue_4 TxQueue ( .Clk_r(Clk_r), .Rst_n(Rst_n), .Packet_In(
        Packet_From_Core), .Read_Ack(TxQueue_Read), .Write_Ack(TxQueue_Write), 
        .Packet_Out(TxData), .Empty(TxQueue_Empty), .Full(TxQueue_Full) );
  Packet_Queue_3 RxQueue ( .Clk_r(Clk_r), .Rst_n(Rst_n), .Packet_In(RxData), 
        .Read_Ack(RxQueue_Read), .Write_Ack(RxQueue_Write), .Packet_Out(
        Packet_To_Core), .Empty(RxQueue_Empty), .Full(RxQueue_Full) );
  FD2QM1P Core_Rcv_Ready_reg ( .D(N9), .CP(Clk_r), .CD(Rst_n), .Q(
        Core_Rcv_Ready) );
  FD2QM1P TxQueue_Read_reg ( .D(N16), .CP(Clk_r), .CD(Rst_n), .Q(TxQueue_Read)
         );
  FD4QM1P RxQueue_Write_reg ( .D(n7), .CP(Clk_r), .SD(Rst_n), .Q(n6) );
  FD4QM1P TxData_Valid_reg ( .D(n9), .CP(Clk_r), .SD(Rst_n), .Q(n8) );
  N1M2P U3 ( .A(n6), .Z(RxQueue_Write) );
  OA21M1P U4 ( .A(Core_Rcv_Ready), .B(n5), .C(n6), .Z(N9) );
  NR2M1P U5 ( .A(n8), .B(Tx_Ready), .Z(N16) );
  NR2M1P U6 ( .A(RxData_Valid), .B(RxQueue_Full), .Z(n5) );
  N1M1P U7 ( .A(n8), .Z(TxData_Valid) );
  ND3M1P U8 ( .A(n6), .B(Core_Rcv_Ready), .C(RxData_Valid), .Z(n7) );
  AO21CNM1P U9 ( .A(n8), .B(TxQueue_Empty), .C(Tx_Ready), .Z(n9) );
endmodule


module Packet_Queue_5 ( Clk_r, Rst_n, Packet_In, Read_Ack, Write_Ack, 
        Packet_Out, Empty, Full );
  input [31:0] Packet_In;
  output [31:0] Packet_Out;
  input Clk_r, Rst_n, Read_Ack, Write_Ack;
  output Empty, Full;
  wire   \Queue[4][31] , \Queue[4][30] , \Queue[4][29] , \Queue[4][28] ,
         \Queue[4][27] , \Queue[4][26] , \Queue[4][25] , \Queue[4][24] ,
         \Queue[4][23] , \Queue[4][22] , \Queue[4][21] , \Queue[4][20] ,
         \Queue[4][19] , \Queue[4][18] , \Queue[4][17] , \Queue[4][16] ,
         \Queue[4][15] , \Queue[4][14] , \Queue[4][13] , \Queue[4][12] ,
         \Queue[4][11] , \Queue[4][10] , \Queue[4][9] , \Queue[4][8] ,
         \Queue[4][7] , \Queue[4][6] , \Queue[4][5] , \Queue[4][4] ,
         \Queue[4][3] , \Queue[4][2] , \Queue[4][1] , \Queue[4][0] ,
         \Queue[3][31] , \Queue[3][30] , \Queue[3][29] , \Queue[3][28] ,
         \Queue[3][27] , \Queue[3][26] , \Queue[3][25] , \Queue[3][24] ,
         \Queue[3][23] , \Queue[3][22] , \Queue[3][21] , \Queue[3][20] ,
         \Queue[3][19] , \Queue[3][18] , \Queue[3][17] , \Queue[3][16] ,
         \Queue[3][15] , \Queue[3][14] , \Queue[3][13] , \Queue[3][12] ,
         \Queue[3][11] , \Queue[3][10] , \Queue[3][9] , \Queue[3][8] ,
         \Queue[3][7] , \Queue[3][6] , \Queue[3][5] , \Queue[3][4] ,
         \Queue[3][3] , \Queue[3][2] , \Queue[3][1] , \Queue[3][0] ,
         \Queue[2][31] , \Queue[2][30] , \Queue[2][29] , \Queue[2][28] ,
         \Queue[2][27] , \Queue[2][26] , \Queue[2][25] , \Queue[2][24] ,
         \Queue[2][23] , \Queue[2][22] , \Queue[2][21] , \Queue[2][20] ,
         \Queue[2][19] , \Queue[2][18] , \Queue[2][17] , \Queue[2][16] ,
         \Queue[2][15] , \Queue[2][14] , \Queue[2][13] , \Queue[2][12] ,
         \Queue[2][11] , \Queue[2][10] , \Queue[2][9] , \Queue[2][8] ,
         \Queue[2][7] , \Queue[2][6] , \Queue[2][5] , \Queue[2][4] ,
         \Queue[2][3] , \Queue[2][2] , \Queue[2][1] , \Queue[2][0] ,
         \Queue[1][31] , \Queue[1][30] , \Queue[1][29] , \Queue[1][28] ,
         \Queue[1][27] , \Queue[1][26] , \Queue[1][25] , \Queue[1][24] ,
         \Queue[1][23] , \Queue[1][22] , \Queue[1][21] , \Queue[1][20] ,
         \Queue[1][19] , \Queue[1][18] , \Queue[1][17] , \Queue[1][16] ,
         \Queue[1][15] , \Queue[1][14] , \Queue[1][13] , \Queue[1][12] ,
         \Queue[1][11] , \Queue[1][10] , \Queue[1][9] , \Queue[1][8] ,
         \Queue[1][7] , \Queue[1][6] , \Queue[1][5] , \Queue[1][4] ,
         \Queue[1][3] , \Queue[1][2] , \Queue[1][1] , \Queue[1][0] , n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541;
  wire   [2:0] Count;

  FDN2QM1P \Count_reg[0]  ( .D(n376), .CPN(Clk_r), .CD(Rst_n), .Q(Count[0]) );
  FDN2QM1P \Count_reg[1]  ( .D(n377), .CPN(Clk_r), .CD(Rst_n), .Q(Count[1]) );
  FDN2QM1P \Count_reg[2]  ( .D(n378), .CPN(Clk_r), .CD(Rst_n), .Q(Count[2]) );
  FDN1QM1P \Queue_reg[4][30]  ( .D(n410), .CPN(Clk_r), .Q(\Queue[4][30] ) );
  FDN1QM1P \Queue_reg[3][30]  ( .D(n538), .CPN(Clk_r), .Q(\Queue[3][30] ) );
  FDN1QM1P \Queue_reg[2][30]  ( .D(n506), .CPN(Clk_r), .Q(\Queue[2][30] ) );
  FDN1QM1P \Queue_reg[4][29]  ( .D(n409), .CPN(Clk_r), .Q(\Queue[4][29] ) );
  FDN1QM1P \Queue_reg[3][29]  ( .D(n537), .CPN(Clk_r), .Q(\Queue[3][29] ) );
  FDN1QM1P \Queue_reg[2][29]  ( .D(n505), .CPN(Clk_r), .Q(\Queue[2][29] ) );
  FDN1QM1P \Queue_reg[4][28]  ( .D(n408), .CPN(Clk_r), .Q(\Queue[4][28] ) );
  FDN1QM1P \Queue_reg[3][28]  ( .D(n536), .CPN(Clk_r), .Q(\Queue[3][28] ) );
  FDN1QM1P \Queue_reg[2][28]  ( .D(n504), .CPN(Clk_r), .Q(\Queue[2][28] ) );
  FDN1QM1P \Queue_reg[4][27]  ( .D(n407), .CPN(Clk_r), .Q(\Queue[4][27] ) );
  FDN1QM1P \Queue_reg[3][27]  ( .D(n535), .CPN(Clk_r), .Q(\Queue[3][27] ) );
  FDN1QM1P \Queue_reg[2][27]  ( .D(n503), .CPN(Clk_r), .Q(\Queue[2][27] ) );
  FDN1QM1P \Queue_reg[4][26]  ( .D(n406), .CPN(Clk_r), .Q(\Queue[4][26] ) );
  FDN1QM1P \Queue_reg[3][26]  ( .D(n534), .CPN(Clk_r), .Q(\Queue[3][26] ) );
  FDN1QM1P \Queue_reg[2][26]  ( .D(n502), .CPN(Clk_r), .Q(\Queue[2][26] ) );
  FDN1QM1P \Queue_reg[4][25]  ( .D(n405), .CPN(Clk_r), .Q(\Queue[4][25] ) );
  FDN1QM1P \Queue_reg[3][25]  ( .D(n533), .CPN(Clk_r), .Q(\Queue[3][25] ) );
  FDN1QM1P \Queue_reg[2][25]  ( .D(n501), .CPN(Clk_r), .Q(\Queue[2][25] ) );
  FDN1QM1P \Queue_reg[4][24]  ( .D(n404), .CPN(Clk_r), .Q(\Queue[4][24] ) );
  FDN1QM1P \Queue_reg[3][24]  ( .D(n532), .CPN(Clk_r), .Q(\Queue[3][24] ) );
  FDN1QM1P \Queue_reg[2][24]  ( .D(n500), .CPN(Clk_r), .Q(\Queue[2][24] ) );
  FDN1QM1P \Queue_reg[4][23]  ( .D(n403), .CPN(Clk_r), .Q(\Queue[4][23] ) );
  FDN1QM1P \Queue_reg[3][23]  ( .D(n531), .CPN(Clk_r), .Q(\Queue[3][23] ) );
  FDN1QM1P \Queue_reg[2][23]  ( .D(n499), .CPN(Clk_r), .Q(\Queue[2][23] ) );
  FDN1QM1P \Queue_reg[4][22]  ( .D(n402), .CPN(Clk_r), .Q(\Queue[4][22] ) );
  FDN1QM1P \Queue_reg[3][22]  ( .D(n530), .CPN(Clk_r), .Q(\Queue[3][22] ) );
  FDN1QM1P \Queue_reg[2][22]  ( .D(n498), .CPN(Clk_r), .Q(\Queue[2][22] ) );
  FDN1QM1P \Queue_reg[4][21]  ( .D(n401), .CPN(Clk_r), .Q(\Queue[4][21] ) );
  FDN1QM1P \Queue_reg[3][21]  ( .D(n529), .CPN(Clk_r), .Q(\Queue[3][21] ) );
  FDN1QM1P \Queue_reg[2][21]  ( .D(n497), .CPN(Clk_r), .Q(\Queue[2][21] ) );
  FDN1QM1P \Queue_reg[4][20]  ( .D(n400), .CPN(Clk_r), .Q(\Queue[4][20] ) );
  FDN1QM1P \Queue_reg[3][20]  ( .D(n528), .CPN(Clk_r), .Q(\Queue[3][20] ) );
  FDN1QM1P \Queue_reg[2][20]  ( .D(n496), .CPN(Clk_r), .Q(\Queue[2][20] ) );
  FDN1QM1P \Queue_reg[4][19]  ( .D(n399), .CPN(Clk_r), .Q(\Queue[4][19] ) );
  FDN1QM1P \Queue_reg[3][19]  ( .D(n527), .CPN(Clk_r), .Q(\Queue[3][19] ) );
  FDN1QM1P \Queue_reg[2][19]  ( .D(n495), .CPN(Clk_r), .Q(\Queue[2][19] ) );
  FDN1QM1P \Queue_reg[4][18]  ( .D(n398), .CPN(Clk_r), .Q(\Queue[4][18] ) );
  FDN1QM1P \Queue_reg[3][18]  ( .D(n526), .CPN(Clk_r), .Q(\Queue[3][18] ) );
  FDN1QM1P \Queue_reg[2][18]  ( .D(n494), .CPN(Clk_r), .Q(\Queue[2][18] ) );
  FDN1QM1P \Queue_reg[4][17]  ( .D(n397), .CPN(Clk_r), .Q(\Queue[4][17] ) );
  FDN1QM1P \Queue_reg[3][17]  ( .D(n525), .CPN(Clk_r), .Q(\Queue[3][17] ) );
  FDN1QM1P \Queue_reg[2][17]  ( .D(n493), .CPN(Clk_r), .Q(\Queue[2][17] ) );
  FDN1QM1P \Queue_reg[4][16]  ( .D(n396), .CPN(Clk_r), .Q(\Queue[4][16] ) );
  FDN1QM1P \Queue_reg[3][16]  ( .D(n524), .CPN(Clk_r), .Q(\Queue[3][16] ) );
  FDN1QM1P \Queue_reg[2][16]  ( .D(n492), .CPN(Clk_r), .Q(\Queue[2][16] ) );
  FDN1QM1P \Queue_reg[4][15]  ( .D(n395), .CPN(Clk_r), .Q(\Queue[4][15] ) );
  FDN1QM1P \Queue_reg[3][15]  ( .D(n523), .CPN(Clk_r), .Q(\Queue[3][15] ) );
  FDN1QM1P \Queue_reg[2][15]  ( .D(n491), .CPN(Clk_r), .Q(\Queue[2][15] ) );
  FDN1QM1P \Queue_reg[4][14]  ( .D(n394), .CPN(Clk_r), .Q(\Queue[4][14] ) );
  FDN1QM1P \Queue_reg[3][14]  ( .D(n522), .CPN(Clk_r), .Q(\Queue[3][14] ) );
  FDN1QM1P \Queue_reg[2][14]  ( .D(n490), .CPN(Clk_r), .Q(\Queue[2][14] ) );
  FDN1QM1P \Queue_reg[4][13]  ( .D(n393), .CPN(Clk_r), .Q(\Queue[4][13] ) );
  FDN1QM1P \Queue_reg[3][13]  ( .D(n521), .CPN(Clk_r), .Q(\Queue[3][13] ) );
  FDN1QM1P \Queue_reg[2][13]  ( .D(n489), .CPN(Clk_r), .Q(\Queue[2][13] ) );
  FDN1QM1P \Queue_reg[4][12]  ( .D(n392), .CPN(Clk_r), .Q(\Queue[4][12] ) );
  FDN1QM1P \Queue_reg[3][12]  ( .D(n520), .CPN(Clk_r), .Q(\Queue[3][12] ) );
  FDN1QM1P \Queue_reg[2][12]  ( .D(n488), .CPN(Clk_r), .Q(\Queue[2][12] ) );
  FDN1QM1P \Queue_reg[4][11]  ( .D(n391), .CPN(Clk_r), .Q(\Queue[4][11] ) );
  FDN1QM1P \Queue_reg[3][11]  ( .D(n519), .CPN(Clk_r), .Q(\Queue[3][11] ) );
  FDN1QM1P \Queue_reg[2][11]  ( .D(n487), .CPN(Clk_r), .Q(\Queue[2][11] ) );
  FDN1QM1P \Queue_reg[4][10]  ( .D(n390), .CPN(Clk_r), .Q(\Queue[4][10] ) );
  FDN1QM1P \Queue_reg[3][10]  ( .D(n518), .CPN(Clk_r), .Q(\Queue[3][10] ) );
  FDN1QM1P \Queue_reg[2][10]  ( .D(n486), .CPN(Clk_r), .Q(\Queue[2][10] ) );
  FDN1QM1P \Queue_reg[4][9]  ( .D(n389), .CPN(Clk_r), .Q(\Queue[4][9] ) );
  FDN1QM1P \Queue_reg[3][9]  ( .D(n517), .CPN(Clk_r), .Q(\Queue[3][9] ) );
  FDN1QM1P \Queue_reg[2][9]  ( .D(n485), .CPN(Clk_r), .Q(\Queue[2][9] ) );
  FDN1QM1P \Queue_reg[4][8]  ( .D(n388), .CPN(Clk_r), .Q(\Queue[4][8] ) );
  FDN1QM1P \Queue_reg[3][8]  ( .D(n516), .CPN(Clk_r), .Q(\Queue[3][8] ) );
  FDN1QM1P \Queue_reg[2][8]  ( .D(n484), .CPN(Clk_r), .Q(\Queue[2][8] ) );
  FDN1QM1P \Queue_reg[4][7]  ( .D(n387), .CPN(Clk_r), .Q(\Queue[4][7] ) );
  FDN1QM1P \Queue_reg[3][7]  ( .D(n515), .CPN(Clk_r), .Q(\Queue[3][7] ) );
  FDN1QM1P \Queue_reg[2][7]  ( .D(n483), .CPN(Clk_r), .Q(\Queue[2][7] ) );
  FDN1QM1P \Queue_reg[4][6]  ( .D(n386), .CPN(Clk_r), .Q(\Queue[4][6] ) );
  FDN1QM1P \Queue_reg[3][6]  ( .D(n514), .CPN(Clk_r), .Q(\Queue[3][6] ) );
  FDN1QM1P \Queue_reg[2][6]  ( .D(n482), .CPN(Clk_r), .Q(\Queue[2][6] ) );
  FDN1QM1P \Queue_reg[4][5]  ( .D(n385), .CPN(Clk_r), .Q(\Queue[4][5] ) );
  FDN1QM1P \Queue_reg[3][5]  ( .D(n513), .CPN(Clk_r), .Q(\Queue[3][5] ) );
  FDN1QM1P \Queue_reg[2][5]  ( .D(n481), .CPN(Clk_r), .Q(\Queue[2][5] ) );
  FDN1QM1P \Queue_reg[4][4]  ( .D(n384), .CPN(Clk_r), .Q(\Queue[4][4] ) );
  FDN1QM1P \Queue_reg[3][4]  ( .D(n512), .CPN(Clk_r), .Q(\Queue[3][4] ) );
  FDN1QM1P \Queue_reg[2][4]  ( .D(n480), .CPN(Clk_r), .Q(\Queue[2][4] ) );
  FDN1QM1P \Queue_reg[4][3]  ( .D(n383), .CPN(Clk_r), .Q(\Queue[4][3] ) );
  FDN1QM1P \Queue_reg[3][3]  ( .D(n511), .CPN(Clk_r), .Q(\Queue[3][3] ) );
  FDN1QM1P \Queue_reg[2][3]  ( .D(n479), .CPN(Clk_r), .Q(\Queue[2][3] ) );
  FDN1QM1P \Queue_reg[4][2]  ( .D(n382), .CPN(Clk_r), .Q(\Queue[4][2] ) );
  FDN1QM1P \Queue_reg[3][2]  ( .D(n510), .CPN(Clk_r), .Q(\Queue[3][2] ) );
  FDN1QM1P \Queue_reg[2][2]  ( .D(n478), .CPN(Clk_r), .Q(\Queue[2][2] ) );
  FDN1QM1P \Queue_reg[4][1]  ( .D(n381), .CPN(Clk_r), .Q(\Queue[4][1] ) );
  FDN1QM1P \Queue_reg[3][1]  ( .D(n509), .CPN(Clk_r), .Q(\Queue[3][1] ) );
  FDN1QM1P \Queue_reg[2][1]  ( .D(n477), .CPN(Clk_r), .Q(\Queue[2][1] ) );
  FDN1QM1P \Queue_reg[4][0]  ( .D(n380), .CPN(Clk_r), .Q(\Queue[4][0] ) );
  FDN1QM1P \Queue_reg[3][0]  ( .D(n508), .CPN(Clk_r), .Q(\Queue[3][0] ) );
  FDN1QM1P \Queue_reg[2][0]  ( .D(n476), .CPN(Clk_r), .Q(\Queue[2][0] ) );
  FDN1QM1P \Queue_reg[4][31]  ( .D(n379), .CPN(Clk_r), .Q(\Queue[4][31] ) );
  FDN1QM1P \Queue_reg[3][31]  ( .D(n539), .CPN(Clk_r), .Q(\Queue[3][31] ) );
  FDN1QM1P \Queue_reg[2][31]  ( .D(n507), .CPN(Clk_r), .Q(\Queue[2][31] ) );
  FDN2QM1P Full_reg ( .D(n411), .CPN(Clk_r), .CD(Rst_n), .Q(Full) );
  FDN1QM1P \Queue_reg[1][31]  ( .D(n443), .CPN(Clk_r), .Q(\Queue[1][31] ) );
  FDN1QM1P \Queue_reg[0][31]  ( .D(n475), .CPN(Clk_r), .Q(Packet_Out[31]) );
  FDN1QM1P \Queue_reg[1][30]  ( .D(n442), .CPN(Clk_r), .Q(\Queue[1][30] ) );
  FDN1QM1P \Queue_reg[0][30]  ( .D(n474), .CPN(Clk_r), .Q(Packet_Out[30]) );
  FDN1QM1P \Queue_reg[1][29]  ( .D(n441), .CPN(Clk_r), .Q(\Queue[1][29] ) );
  FDN1QM1P \Queue_reg[0][29]  ( .D(n473), .CPN(Clk_r), .Q(Packet_Out[29]) );
  FDN1QM1P \Queue_reg[1][28]  ( .D(n440), .CPN(Clk_r), .Q(\Queue[1][28] ) );
  FDN1QM1P \Queue_reg[0][28]  ( .D(n472), .CPN(Clk_r), .Q(Packet_Out[28]) );
  FDN1QM1P \Queue_reg[1][27]  ( .D(n439), .CPN(Clk_r), .Q(\Queue[1][27] ) );
  FDN1QM1P \Queue_reg[0][27]  ( .D(n471), .CPN(Clk_r), .Q(Packet_Out[27]) );
  FDN1QM1P \Queue_reg[1][26]  ( .D(n438), .CPN(Clk_r), .Q(\Queue[1][26] ) );
  FDN1QM1P \Queue_reg[0][26]  ( .D(n470), .CPN(Clk_r), .Q(Packet_Out[26]) );
  FDN1QM1P \Queue_reg[1][25]  ( .D(n437), .CPN(Clk_r), .Q(\Queue[1][25] ) );
  FDN1QM1P \Queue_reg[0][25]  ( .D(n469), .CPN(Clk_r), .Q(Packet_Out[25]) );
  FDN1QM1P \Queue_reg[1][24]  ( .D(n436), .CPN(Clk_r), .Q(\Queue[1][24] ) );
  FDN1QM1P \Queue_reg[0][24]  ( .D(n468), .CPN(Clk_r), .Q(Packet_Out[24]) );
  FDN1QM1P \Queue_reg[1][23]  ( .D(n435), .CPN(Clk_r), .Q(\Queue[1][23] ) );
  FDN1QM1P \Queue_reg[0][23]  ( .D(n467), .CPN(Clk_r), .Q(Packet_Out[23]) );
  FDN1QM1P \Queue_reg[1][22]  ( .D(n434), .CPN(Clk_r), .Q(\Queue[1][22] ) );
  FDN1QM1P \Queue_reg[0][22]  ( .D(n466), .CPN(Clk_r), .Q(Packet_Out[22]) );
  FDN1QM1P \Queue_reg[1][21]  ( .D(n433), .CPN(Clk_r), .Q(\Queue[1][21] ) );
  FDN1QM1P \Queue_reg[0][21]  ( .D(n465), .CPN(Clk_r), .Q(Packet_Out[21]) );
  FDN1QM1P \Queue_reg[1][20]  ( .D(n432), .CPN(Clk_r), .Q(\Queue[1][20] ) );
  FDN1QM1P \Queue_reg[0][20]  ( .D(n464), .CPN(Clk_r), .Q(Packet_Out[20]) );
  FDN1QM1P \Queue_reg[1][19]  ( .D(n431), .CPN(Clk_r), .Q(\Queue[1][19] ) );
  FDN1QM1P \Queue_reg[0][19]  ( .D(n463), .CPN(Clk_r), .Q(Packet_Out[19]) );
  FDN1QM1P \Queue_reg[1][18]  ( .D(n430), .CPN(Clk_r), .Q(\Queue[1][18] ) );
  FDN1QM1P \Queue_reg[0][18]  ( .D(n462), .CPN(Clk_r), .Q(Packet_Out[18]) );
  FDN1QM1P \Queue_reg[1][17]  ( .D(n429), .CPN(Clk_r), .Q(\Queue[1][17] ) );
  FDN1QM1P \Queue_reg[0][17]  ( .D(n461), .CPN(Clk_r), .Q(Packet_Out[17]) );
  FDN1QM1P \Queue_reg[1][16]  ( .D(n428), .CPN(Clk_r), .Q(\Queue[1][16] ) );
  FDN1QM1P \Queue_reg[0][16]  ( .D(n460), .CPN(Clk_r), .Q(Packet_Out[16]) );
  FDN1QM1P \Queue_reg[1][15]  ( .D(n427), .CPN(Clk_r), .Q(\Queue[1][15] ) );
  FDN1QM1P \Queue_reg[0][15]  ( .D(n459), .CPN(Clk_r), .Q(Packet_Out[15]) );
  FDN1QM1P \Queue_reg[1][14]  ( .D(n426), .CPN(Clk_r), .Q(\Queue[1][14] ) );
  FDN1QM1P \Queue_reg[0][14]  ( .D(n458), .CPN(Clk_r), .Q(Packet_Out[14]) );
  FDN1QM1P \Queue_reg[1][13]  ( .D(n425), .CPN(Clk_r), .Q(\Queue[1][13] ) );
  FDN1QM1P \Queue_reg[0][13]  ( .D(n457), .CPN(Clk_r), .Q(Packet_Out[13]) );
  FDN1QM1P \Queue_reg[1][12]  ( .D(n424), .CPN(Clk_r), .Q(\Queue[1][12] ) );
  FDN1QM1P \Queue_reg[0][12]  ( .D(n456), .CPN(Clk_r), .Q(Packet_Out[12]) );
  FDN1QM1P \Queue_reg[1][11]  ( .D(n423), .CPN(Clk_r), .Q(\Queue[1][11] ) );
  FDN1QM1P \Queue_reg[0][11]  ( .D(n455), .CPN(Clk_r), .Q(Packet_Out[11]) );
  FDN1QM1P \Queue_reg[1][10]  ( .D(n422), .CPN(Clk_r), .Q(\Queue[1][10] ) );
  FDN1QM1P \Queue_reg[0][10]  ( .D(n454), .CPN(Clk_r), .Q(Packet_Out[10]) );
  FDN1QM1P \Queue_reg[1][9]  ( .D(n421), .CPN(Clk_r), .Q(\Queue[1][9] ) );
  FDN1QM1P \Queue_reg[0][9]  ( .D(n453), .CPN(Clk_r), .Q(Packet_Out[9]) );
  FDN1QM1P \Queue_reg[1][8]  ( .D(n420), .CPN(Clk_r), .Q(\Queue[1][8] ) );
  FDN1QM1P \Queue_reg[0][8]  ( .D(n452), .CPN(Clk_r), .Q(Packet_Out[8]) );
  FDN1QM1P \Queue_reg[1][7]  ( .D(n419), .CPN(Clk_r), .Q(\Queue[1][7] ) );
  FDN1QM1P \Queue_reg[0][7]  ( .D(n451), .CPN(Clk_r), .Q(Packet_Out[7]) );
  FDN1QM1P \Queue_reg[1][6]  ( .D(n418), .CPN(Clk_r), .Q(\Queue[1][6] ) );
  FDN1QM1P \Queue_reg[0][6]  ( .D(n450), .CPN(Clk_r), .Q(Packet_Out[6]) );
  FDN1QM1P \Queue_reg[1][5]  ( .D(n417), .CPN(Clk_r), .Q(\Queue[1][5] ) );
  FDN1QM1P \Queue_reg[0][5]  ( .D(n449), .CPN(Clk_r), .Q(Packet_Out[5]) );
  FDN1QM1P \Queue_reg[1][4]  ( .D(n416), .CPN(Clk_r), .Q(\Queue[1][4] ) );
  FDN1QM1P \Queue_reg[0][4]  ( .D(n448), .CPN(Clk_r), .Q(Packet_Out[4]) );
  FDN1QM1P \Queue_reg[1][3]  ( .D(n415), .CPN(Clk_r), .Q(\Queue[1][3] ) );
  FDN1QM1P \Queue_reg[0][3]  ( .D(n447), .CPN(Clk_r), .Q(Packet_Out[3]) );
  FDN1QM1P \Queue_reg[1][2]  ( .D(n414), .CPN(Clk_r), .Q(\Queue[1][2] ) );
  FDN1QM1P \Queue_reg[0][2]  ( .D(n446), .CPN(Clk_r), .Q(Packet_Out[2]) );
  FDN1QM1P \Queue_reg[1][1]  ( .D(n413), .CPN(Clk_r), .Q(\Queue[1][1] ) );
  FDN1QM1P \Queue_reg[0][1]  ( .D(n445), .CPN(Clk_r), .Q(Packet_Out[1]) );
  FDN1QM1P \Queue_reg[1][0]  ( .D(n412), .CPN(Clk_r), .Q(\Queue[1][0] ) );
  FDN1QM1P \Queue_reg[0][0]  ( .D(n444), .CPN(Clk_r), .Q(Packet_Out[0]) );
  FDN2QM1P Empty_reg ( .D(n541), .CPN(Clk_r), .CD(Rst_n), .Q(n540) );
  BUFM2P U3 ( .A(n96), .Z(n8) );
  BUFM1P U4 ( .A(n96), .Z(n9) );
  BUFM1P U5 ( .A(n205), .Z(n11) );
  BUFM2P U6 ( .A(n205), .Z(n10) );
  N1M1P U7 ( .A(Read_Ack), .Z(n136) );
  AOI21M3P U8 ( .A(Write_Ack), .B(n375), .C(n140), .Z(n94) );
  OAI211M4P U9 ( .A(n139), .B(n136), .C(Write_Ack), .D(n97), .Z(n134) );
  OAI211M4P U10 ( .A(n141), .B(n136), .C(Write_Ack), .D(n135), .Z(n207) );
  AOI21M3P U11 ( .A(Write_Ack), .B(n99), .C(n140), .Z(n56) );
  AOI21M3P U12 ( .A(Write_Ack), .B(n141), .C(n140), .Z(n204) );
  AOI21M3P U13 ( .A(Write_Ack), .B(n139), .C(n140), .Z(n131) );
  OAI211M4P U14 ( .A(n99), .B(n138), .C(Rst_n), .D(n137), .Z(n132) );
  NR2I1M8P U15 ( .A(n60), .B(n20), .Z(n19) );
  OAI211M4P U16 ( .A(n99), .B(n136), .C(Write_Ack), .D(n23), .Z(n58) );
  ND2M1P U17 ( .A(n17), .B(Rst_n), .Z(n60) );
  NR2M2P U18 ( .A(Read_Ack), .B(n98), .Z(n17) );
  NR3M1P U19 ( .A(n22), .B(Count[2]), .C(Count[1]), .Z(n375) );
  NR3M1P U20 ( .A(Count[2]), .B(n22), .C(n21), .Z(n139) );
  NR3M1P U21 ( .A(Count[0]), .B(Count[2]), .C(n21), .Z(n99) );
  NR3M1P U22 ( .A(Count[0]), .B(Count[1]), .C(n18), .Z(n141) );
  N1M1P U23 ( .A(Count[0]), .Z(n22) );
  N1M1P U24 ( .A(Count[1]), .Z(n21) );
  N1M1P U25 ( .A(Count[2]), .Z(n18) );
  ND2M2P U26 ( .A(Read_Ack), .B(Rst_n), .Z(n140) );
  BUFM2P U27 ( .A(n55), .Z(n3) );
  BUFM2P U28 ( .A(n55), .Z(n5) );
  BUFM2P U29 ( .A(n55), .Z(n4) );
  N1M2P U30 ( .A(n17), .Z(n138) );
  BUFM2P U31 ( .A(n93), .Z(n6) );
  BUFM2P U32 ( .A(n93), .Z(n7) );
  OAI211M1P U33 ( .A(n375), .B(n136), .C(Write_Ack), .D(n61), .Z(n96) );
  N1M2P U34 ( .A(Write_Ack), .Z(n98) );
  OAI211M1P U35 ( .A(n139), .B(n138), .C(Rst_n), .D(n137), .Z(n205) );
  NR2M1P U36 ( .A(n136), .B(Write_Ack), .Z(n374) );
  NR2M1P U37 ( .A(n17), .B(n374), .Z(n373) );
  AOI22CDNM1P U38 ( .A(n373), .B(n22), .C(n373), .D(n22), .Z(n376) );
  N1M1P U39 ( .A(n374), .Z(n16) );
  AOI22M1P U40 ( .A(Count[0]), .B(n138), .C(n16), .D(n22), .Z(n13) );
  AOI22CDNM1P U41 ( .A(Count[1]), .B(n13), .C(n13), .D(Count[1]), .Z(n377) );
  ND3M1P U42 ( .A(n22), .B(n18), .C(n21), .Z(n59) );
  ND2M1P U43 ( .A(Count[1]), .B(Read_Ack), .Z(n12) );
  OAI211M1P U44 ( .A(Count[1]), .B(n138), .C(n13), .D(n12), .Z(n14) );
  AOI22M1P U45 ( .A(n17), .B(n139), .C(Count[2]), .D(n14), .Z(n15) );
  OAI21M1P U46 ( .A(n59), .B(n16), .C(n15), .Z(n378) );
  N1M1P U47 ( .A(n141), .Z(n20) );
  N1M1P U48 ( .A(Packet_In[31]), .Z(n208) );
  AOI22CDNM1P U49 ( .A(n19), .B(n208), .C(\Queue[4][31] ), .D(n19), .Z(n379)
         );
  N1M1P U50 ( .A(Packet_In[0]), .Z(n143) );
  AOI22CDNM1P U51 ( .A(n19), .B(n143), .C(\Queue[4][0] ), .D(n19), .Z(n380) );
  N1M1P U52 ( .A(Packet_In[1]), .Z(n145) );
  AOI22CDNM1P U53 ( .A(n19), .B(n145), .C(\Queue[4][1] ), .D(n19), .Z(n381) );
  N1M1P U54 ( .A(Packet_In[2]), .Z(n147) );
  AOI22CDNM1P U55 ( .A(n19), .B(n147), .C(\Queue[4][2] ), .D(n19), .Z(n382) );
  N1M1P U56 ( .A(Packet_In[3]), .Z(n149) );
  AOI22CDNM1P U57 ( .A(n19), .B(n149), .C(\Queue[4][3] ), .D(n19), .Z(n383) );
  N1M1P U58 ( .A(Packet_In[4]), .Z(n151) );
  AOI22CDNM1P U59 ( .A(n19), .B(n151), .C(\Queue[4][4] ), .D(n19), .Z(n384) );
  N1M1P U60 ( .A(Packet_In[5]), .Z(n153) );
  AOI22CDNM1P U61 ( .A(n19), .B(n153), .C(\Queue[4][5] ), .D(n19), .Z(n385) );
  N1M1P U62 ( .A(Packet_In[6]), .Z(n155) );
  AOI22CDNM1P U63 ( .A(n19), .B(n155), .C(\Queue[4][6] ), .D(n19), .Z(n386) );
  N1M1P U64 ( .A(Packet_In[7]), .Z(n157) );
  AOI22CDNM1P U65 ( .A(n19), .B(n157), .C(\Queue[4][7] ), .D(n19), .Z(n387) );
  N1M1P U66 ( .A(Packet_In[8]), .Z(n159) );
  AOI22CDNM1P U67 ( .A(n19), .B(n159), .C(\Queue[4][8] ), .D(n19), .Z(n388) );
  N1M1P U68 ( .A(Packet_In[9]), .Z(n161) );
  AOI22CDNM1P U69 ( .A(n19), .B(n161), .C(\Queue[4][9] ), .D(n19), .Z(n389) );
  N1M1P U70 ( .A(Packet_In[10]), .Z(n163) );
  AOI22CDNM1P U71 ( .A(n19), .B(n163), .C(\Queue[4][10] ), .D(n19), .Z(n390)
         );
  N1M1P U72 ( .A(Packet_In[11]), .Z(n165) );
  AOI22CDNM1P U73 ( .A(n19), .B(n165), .C(\Queue[4][11] ), .D(n19), .Z(n391)
         );
  N1M1P U74 ( .A(Packet_In[12]), .Z(n167) );
  AOI22CDNM1P U75 ( .A(n19), .B(n167), .C(\Queue[4][12] ), .D(n19), .Z(n392)
         );
  N1M1P U76 ( .A(Packet_In[13]), .Z(n169) );
  AOI22CDNM1P U77 ( .A(n19), .B(n169), .C(\Queue[4][13] ), .D(n19), .Z(n393)
         );
  N1M1P U78 ( .A(Packet_In[14]), .Z(n171) );
  AOI22CDNM1P U79 ( .A(n19), .B(n171), .C(\Queue[4][14] ), .D(n19), .Z(n394)
         );
  N1M1P U80 ( .A(Packet_In[15]), .Z(n173) );
  AOI22CDNM1P U81 ( .A(n19), .B(n173), .C(\Queue[4][15] ), .D(n19), .Z(n395)
         );
  N1M1P U82 ( .A(Packet_In[16]), .Z(n175) );
  AOI22CDNM1P U83 ( .A(n19), .B(n175), .C(\Queue[4][16] ), .D(n19), .Z(n396)
         );
  N1M1P U84 ( .A(Packet_In[17]), .Z(n177) );
  AOI22CDNM1P U85 ( .A(n19), .B(n177), .C(\Queue[4][17] ), .D(n19), .Z(n397)
         );
  N1M1P U86 ( .A(Packet_In[18]), .Z(n179) );
  AOI22CDNM1P U87 ( .A(n19), .B(n179), .C(\Queue[4][18] ), .D(n19), .Z(n398)
         );
  N1M1P U88 ( .A(Packet_In[19]), .Z(n181) );
  AOI22CDNM1P U89 ( .A(n19), .B(n181), .C(\Queue[4][19] ), .D(n19), .Z(n399)
         );
  N1M1P U90 ( .A(Packet_In[20]), .Z(n183) );
  AOI22CDNM1P U91 ( .A(n19), .B(n183), .C(\Queue[4][20] ), .D(n19), .Z(n400)
         );
  N1M1P U92 ( .A(Packet_In[21]), .Z(n185) );
  AOI22CDNM1P U93 ( .A(n19), .B(n185), .C(\Queue[4][21] ), .D(n19), .Z(n401)
         );
  N1M1P U94 ( .A(Packet_In[22]), .Z(n187) );
  AOI22CDNM1P U95 ( .A(n19), .B(n187), .C(\Queue[4][22] ), .D(n19), .Z(n402)
         );
  N1M1P U96 ( .A(Packet_In[23]), .Z(n189) );
  AOI22CDNM1P U97 ( .A(n19), .B(n189), .C(\Queue[4][23] ), .D(n19), .Z(n403)
         );
  N1M1P U98 ( .A(Packet_In[24]), .Z(n191) );
  AOI22CDNM1P U99 ( .A(n19), .B(n191), .C(\Queue[4][24] ), .D(n19), .Z(n404)
         );
  N1M1P U100 ( .A(Packet_In[25]), .Z(n193) );
  AOI22CDNM1P U101 ( .A(n19), .B(n193), .C(\Queue[4][25] ), .D(n19), .Z(n405)
         );
  N1M1P U102 ( .A(Packet_In[26]), .Z(n195) );
  AOI22CDNM1P U103 ( .A(n19), .B(n195), .C(\Queue[4][26] ), .D(n19), .Z(n406)
         );
  N1M1P U104 ( .A(Packet_In[27]), .Z(n197) );
  AOI22CDNM1P U105 ( .A(n19), .B(n197), .C(\Queue[4][27] ), .D(n19), .Z(n407)
         );
  N1M1P U106 ( .A(Packet_In[28]), .Z(n199) );
  AOI22CDNM1P U107 ( .A(n19), .B(n199), .C(\Queue[4][28] ), .D(n19), .Z(n408)
         );
  N1M1P U108 ( .A(Packet_In[29]), .Z(n201) );
  AOI22CDNM1P U109 ( .A(n19), .B(n201), .C(\Queue[4][29] ), .D(n19), .Z(n409)
         );
  N1M1P U110 ( .A(Packet_In[30]), .Z(n203) );
  AOI22CDNM1P U111 ( .A(n19), .B(n203), .C(\Queue[4][30] ), .D(n19), .Z(n410)
         );
  OAI22CDNM1P U112 ( .A(n138), .B(n20), .C(n373), .D(Full), .Z(n411) );
  OA21M1P U113 ( .A(n138), .B(n375), .C(Rst_n), .Z(n23) );
  OAI21M1P U114 ( .A(Write_Ack), .B(Read_Ack), .C(n23), .Z(n55) );
  AOI22M1P U115 ( .A(\Queue[2][0] ), .B(n56), .C(\Queue[1][0] ), .D(n3), .Z(
        n24) );
  OAI21M1P U116 ( .A(n143), .B(n58), .C(n24), .Z(n412) );
  AOI22M1P U117 ( .A(n56), .B(\Queue[2][1] ), .C(\Queue[1][1] ), .D(n3), .Z(
        n25) );
  OAI21M1P U118 ( .A(n58), .B(n145), .C(n25), .Z(n413) );
  AOI22M1P U119 ( .A(n56), .B(\Queue[2][2] ), .C(\Queue[1][2] ), .D(n3), .Z(
        n26) );
  OAI21M1P U120 ( .A(n58), .B(n147), .C(n26), .Z(n414) );
  AOI22M1P U121 ( .A(n56), .B(\Queue[2][3] ), .C(\Queue[1][3] ), .D(n3), .Z(
        n27) );
  OAI21M1P U122 ( .A(n58), .B(n149), .C(n27), .Z(n415) );
  AOI22M1P U123 ( .A(n56), .B(\Queue[2][4] ), .C(\Queue[1][4] ), .D(n3), .Z(
        n28) );
  OAI21M1P U124 ( .A(n58), .B(n151), .C(n28), .Z(n416) );
  AOI22M1P U125 ( .A(n56), .B(\Queue[2][5] ), .C(\Queue[1][5] ), .D(n3), .Z(
        n29) );
  OAI21M1P U126 ( .A(n58), .B(n153), .C(n29), .Z(n417) );
  AOI22M1P U127 ( .A(n56), .B(\Queue[2][6] ), .C(\Queue[1][6] ), .D(n3), .Z(
        n30) );
  OAI21M1P U128 ( .A(n58), .B(n155), .C(n30), .Z(n418) );
  AOI22M1P U129 ( .A(n56), .B(\Queue[2][7] ), .C(\Queue[1][7] ), .D(n3), .Z(
        n31) );
  OAI21M1P U130 ( .A(n58), .B(n157), .C(n31), .Z(n419) );
  AOI22M1P U131 ( .A(n56), .B(\Queue[2][8] ), .C(\Queue[1][8] ), .D(n3), .Z(
        n32) );
  OAI21M1P U132 ( .A(n58), .B(n159), .C(n32), .Z(n420) );
  AOI22M1P U133 ( .A(n56), .B(\Queue[2][9] ), .C(\Queue[1][9] ), .D(n4), .Z(
        n33) );
  OAI21M1P U134 ( .A(n58), .B(n161), .C(n33), .Z(n421) );
  AOI22M1P U135 ( .A(n56), .B(\Queue[2][10] ), .C(\Queue[1][10] ), .D(n4), .Z(
        n34) );
  OAI21M1P U136 ( .A(n58), .B(n163), .C(n34), .Z(n422) );
  AOI22M1P U137 ( .A(n56), .B(\Queue[2][11] ), .C(\Queue[1][11] ), .D(n4), .Z(
        n35) );
  OAI21M1P U138 ( .A(n58), .B(n165), .C(n35), .Z(n423) );
  AOI22M1P U139 ( .A(n56), .B(\Queue[2][12] ), .C(\Queue[1][12] ), .D(n4), .Z(
        n36) );
  OAI21M1P U140 ( .A(n58), .B(n167), .C(n36), .Z(n424) );
  AOI22M1P U141 ( .A(n56), .B(\Queue[2][13] ), .C(\Queue[1][13] ), .D(n4), .Z(
        n37) );
  OAI21M1P U142 ( .A(n58), .B(n169), .C(n37), .Z(n425) );
  AOI22M1P U143 ( .A(n56), .B(\Queue[2][14] ), .C(\Queue[1][14] ), .D(n4), .Z(
        n38) );
  OAI21M1P U144 ( .A(n58), .B(n171), .C(n38), .Z(n426) );
  AOI22M1P U145 ( .A(n56), .B(\Queue[2][15] ), .C(\Queue[1][15] ), .D(n4), .Z(
        n39) );
  OAI21M1P U146 ( .A(n58), .B(n173), .C(n39), .Z(n427) );
  AOI22M1P U147 ( .A(n56), .B(\Queue[2][16] ), .C(\Queue[1][16] ), .D(n4), .Z(
        n40) );
  OAI21M1P U148 ( .A(n58), .B(n175), .C(n40), .Z(n428) );
  AOI22M1P U149 ( .A(n56), .B(\Queue[2][17] ), .C(\Queue[1][17] ), .D(n4), .Z(
        n41) );
  OAI21M1P U150 ( .A(n58), .B(n177), .C(n41), .Z(n429) );
  AOI22M1P U151 ( .A(n56), .B(\Queue[2][18] ), .C(\Queue[1][18] ), .D(n5), .Z(
        n42) );
  OAI21M1P U152 ( .A(n58), .B(n179), .C(n42), .Z(n430) );
  AOI22M1P U153 ( .A(n56), .B(\Queue[2][19] ), .C(\Queue[1][19] ), .D(n5), .Z(
        n43) );
  OAI21M1P U154 ( .A(n58), .B(n181), .C(n43), .Z(n431) );
  AOI22M1P U155 ( .A(n56), .B(\Queue[2][20] ), .C(\Queue[1][20] ), .D(n5), .Z(
        n44) );
  OAI21M1P U156 ( .A(n58), .B(n183), .C(n44), .Z(n432) );
  AOI22M1P U157 ( .A(n56), .B(\Queue[2][21] ), .C(\Queue[1][21] ), .D(n5), .Z(
        n45) );
  OAI21M1P U158 ( .A(n58), .B(n185), .C(n45), .Z(n433) );
  AOI22M1P U159 ( .A(n56), .B(\Queue[2][22] ), .C(\Queue[1][22] ), .D(n5), .Z(
        n46) );
  OAI21M1P U160 ( .A(n58), .B(n187), .C(n46), .Z(n434) );
  AOI22M1P U161 ( .A(n56), .B(\Queue[2][23] ), .C(\Queue[1][23] ), .D(n5), .Z(
        n47) );
  OAI21M1P U162 ( .A(n58), .B(n189), .C(n47), .Z(n435) );
  AOI22M1P U163 ( .A(n56), .B(\Queue[2][24] ), .C(\Queue[1][24] ), .D(n5), .Z(
        n48) );
  OAI21M1P U164 ( .A(n58), .B(n191), .C(n48), .Z(n436) );
  AOI22M1P U165 ( .A(n56), .B(\Queue[2][25] ), .C(\Queue[1][25] ), .D(n5), .Z(
        n49) );
  OAI21M1P U166 ( .A(n58), .B(n193), .C(n49), .Z(n437) );
  AOI22M1P U167 ( .A(n56), .B(\Queue[2][26] ), .C(\Queue[1][26] ), .D(n5), .Z(
        n50) );
  OAI21M1P U168 ( .A(n58), .B(n195), .C(n50), .Z(n438) );
  AOI22M1P U169 ( .A(n56), .B(\Queue[2][27] ), .C(\Queue[1][27] ), .D(n4), .Z(
        n51) );
  OAI21M1P U170 ( .A(n58), .B(n197), .C(n51), .Z(n439) );
  AOI22M1P U171 ( .A(n56), .B(\Queue[2][28] ), .C(\Queue[1][28] ), .D(n5), .Z(
        n52) );
  OAI21M1P U172 ( .A(n58), .B(n199), .C(n52), .Z(n440) );
  AOI22M1P U173 ( .A(n56), .B(\Queue[2][29] ), .C(\Queue[1][29] ), .D(n3), .Z(
        n53) );
  OAI21M1P U174 ( .A(n58), .B(n201), .C(n53), .Z(n441) );
  AOI22M1P U175 ( .A(n56), .B(\Queue[2][30] ), .C(\Queue[1][30] ), .D(n4), .Z(
        n54) );
  OAI21M1P U176 ( .A(n58), .B(n203), .C(n54), .Z(n442) );
  AOI22M1P U177 ( .A(n56), .B(\Queue[2][31] ), .C(\Queue[1][31] ), .D(n5), .Z(
        n57) );
  OAI21M1P U178 ( .A(n58), .B(n208), .C(n57), .Z(n443) );
  OAI21M1P U179 ( .A(n60), .B(n59), .C(n140), .Z(n61) );
  N1M1P U180 ( .A(n61), .Z(n93) );
  AOI22M1P U181 ( .A(\Queue[1][0] ), .B(n94), .C(n93), .D(Packet_Out[0]), .Z(
        n62) );
  OAI21M1P U182 ( .A(n143), .B(n8), .C(n62), .Z(n444) );
  AOI22M1P U183 ( .A(\Queue[1][1] ), .B(n94), .C(n93), .D(Packet_Out[1]), .Z(
        n63) );
  OAI21M1P U184 ( .A(n145), .B(n8), .C(n63), .Z(n445) );
  AOI22M1P U185 ( .A(\Queue[1][2] ), .B(n94), .C(n93), .D(Packet_Out[2]), .Z(
        n64) );
  OAI21M1P U186 ( .A(n147), .B(n8), .C(n64), .Z(n446) );
  AOI22M1P U187 ( .A(\Queue[1][3] ), .B(n94), .C(n93), .D(Packet_Out[3]), .Z(
        n65) );
  OAI21M1P U188 ( .A(n149), .B(n8), .C(n65), .Z(n447) );
  AOI22M1P U189 ( .A(\Queue[1][4] ), .B(n94), .C(n93), .D(Packet_Out[4]), .Z(
        n66) );
  OAI21M1P U190 ( .A(n151), .B(n8), .C(n66), .Z(n448) );
  AOI22M1P U191 ( .A(\Queue[1][5] ), .B(n94), .C(n93), .D(Packet_Out[5]), .Z(
        n67) );
  OAI21M1P U192 ( .A(n153), .B(n8), .C(n67), .Z(n449) );
  AOI22M1P U193 ( .A(\Queue[1][6] ), .B(n94), .C(n6), .D(Packet_Out[6]), .Z(
        n68) );
  OAI21M1P U194 ( .A(n155), .B(n8), .C(n68), .Z(n450) );
  AOI22M1P U195 ( .A(\Queue[1][7] ), .B(n94), .C(n7), .D(Packet_Out[7]), .Z(
        n69) );
  OAI21M1P U196 ( .A(n157), .B(n8), .C(n69), .Z(n451) );
  AOI22M1P U197 ( .A(\Queue[1][8] ), .B(n94), .C(n6), .D(Packet_Out[8]), .Z(
        n70) );
  OAI21M1P U198 ( .A(n159), .B(n8), .C(n70), .Z(n452) );
  AOI22M1P U199 ( .A(\Queue[1][9] ), .B(n94), .C(n7), .D(Packet_Out[9]), .Z(
        n71) );
  OAI21M1P U200 ( .A(n161), .B(n8), .C(n71), .Z(n453) );
  AOI22M1P U201 ( .A(\Queue[1][10] ), .B(n94), .C(n6), .D(Packet_Out[10]), .Z(
        n72) );
  OAI21M1P U202 ( .A(n163), .B(n8), .C(n72), .Z(n454) );
  AOI22M1P U203 ( .A(\Queue[1][11] ), .B(n94), .C(n6), .D(Packet_Out[11]), .Z(
        n73) );
  OAI21M1P U204 ( .A(n165), .B(n8), .C(n73), .Z(n455) );
  AOI22M1P U205 ( .A(\Queue[1][12] ), .B(n94), .C(n6), .D(Packet_Out[12]), .Z(
        n74) );
  OAI21M1P U206 ( .A(n167), .B(n8), .C(n74), .Z(n456) );
  AOI22M1P U207 ( .A(\Queue[1][13] ), .B(n94), .C(n6), .D(Packet_Out[13]), .Z(
        n75) );
  OAI21M1P U208 ( .A(n169), .B(n8), .C(n75), .Z(n457) );
  AOI22M1P U209 ( .A(\Queue[1][14] ), .B(n94), .C(n6), .D(Packet_Out[14]), .Z(
        n76) );
  OAI21M1P U210 ( .A(n171), .B(n8), .C(n76), .Z(n458) );
  AOI22M1P U211 ( .A(\Queue[1][15] ), .B(n94), .C(n6), .D(Packet_Out[15]), .Z(
        n77) );
  OAI21M1P U212 ( .A(n173), .B(n8), .C(n77), .Z(n459) );
  AOI22M1P U213 ( .A(\Queue[1][16] ), .B(n94), .C(n6), .D(Packet_Out[16]), .Z(
        n78) );
  OAI21M1P U214 ( .A(n175), .B(n8), .C(n78), .Z(n460) );
  AOI22M1P U215 ( .A(\Queue[1][17] ), .B(n94), .C(n6), .D(Packet_Out[17]), .Z(
        n79) );
  OAI21M1P U216 ( .A(n177), .B(n8), .C(n79), .Z(n461) );
  AOI22M1P U217 ( .A(\Queue[1][18] ), .B(n94), .C(n6), .D(Packet_Out[18]), .Z(
        n80) );
  OAI21M1P U218 ( .A(n179), .B(n8), .C(n80), .Z(n462) );
  AOI22M1P U219 ( .A(\Queue[1][19] ), .B(n94), .C(n6), .D(Packet_Out[19]), .Z(
        n81) );
  OAI21M1P U220 ( .A(n181), .B(n8), .C(n81), .Z(n463) );
  AOI22M1P U221 ( .A(\Queue[1][20] ), .B(n94), .C(n7), .D(Packet_Out[20]), .Z(
        n82) );
  OAI21M1P U222 ( .A(n183), .B(n9), .C(n82), .Z(n464) );
  AOI22M1P U223 ( .A(\Queue[1][21] ), .B(n94), .C(n7), .D(Packet_Out[21]), .Z(
        n83) );
  OAI21M1P U224 ( .A(n185), .B(n9), .C(n83), .Z(n465) );
  AOI22M1P U225 ( .A(\Queue[1][22] ), .B(n94), .C(n7), .D(Packet_Out[22]), .Z(
        n84) );
  OAI21M1P U226 ( .A(n187), .B(n9), .C(n84), .Z(n466) );
  AOI22M1P U227 ( .A(\Queue[1][23] ), .B(n94), .C(n7), .D(Packet_Out[23]), .Z(
        n85) );
  OAI21M1P U228 ( .A(n189), .B(n9), .C(n85), .Z(n467) );
  AOI22M1P U229 ( .A(\Queue[1][24] ), .B(n94), .C(n7), .D(Packet_Out[24]), .Z(
        n86) );
  OAI21M1P U230 ( .A(n191), .B(n9), .C(n86), .Z(n468) );
  AOI22M1P U231 ( .A(\Queue[1][25] ), .B(n94), .C(n7), .D(Packet_Out[25]), .Z(
        n87) );
  OAI21M1P U232 ( .A(n193), .B(n9), .C(n87), .Z(n469) );
  AOI22M1P U233 ( .A(\Queue[1][26] ), .B(n94), .C(n7), .D(Packet_Out[26]), .Z(
        n88) );
  OAI21M1P U234 ( .A(n195), .B(n9), .C(n88), .Z(n470) );
  AOI22M1P U235 ( .A(\Queue[1][27] ), .B(n94), .C(n7), .D(Packet_Out[27]), .Z(
        n89) );
  OAI21M1P U236 ( .A(n197), .B(n9), .C(n89), .Z(n471) );
  AOI22M1P U237 ( .A(\Queue[1][28] ), .B(n94), .C(n7), .D(Packet_Out[28]), .Z(
        n90) );
  OAI21M1P U238 ( .A(n199), .B(n9), .C(n90), .Z(n472) );
  AOI22M1P U239 ( .A(\Queue[1][29] ), .B(n94), .C(n7), .D(Packet_Out[29]), .Z(
        n91) );
  OAI21M1P U240 ( .A(n201), .B(n9), .C(n91), .Z(n473) );
  AOI22M1P U241 ( .A(\Queue[1][30] ), .B(n94), .C(n6), .D(Packet_Out[30]), .Z(
        n92) );
  OAI21M1P U242 ( .A(n203), .B(n8), .C(n92), .Z(n474) );
  AOI22M1P U243 ( .A(\Queue[1][31] ), .B(n94), .C(n7), .D(Packet_Out[31]), .Z(
        n95) );
  OAI21M1P U244 ( .A(n208), .B(n9), .C(n95), .Z(n475) );
  OA21M1P U245 ( .A(n138), .B(n99), .C(Rst_n), .Z(n97) );
  ND2M1P U246 ( .A(n98), .B(n136), .Z(n137) );
  AOI22M1P U247 ( .A(\Queue[2][0] ), .B(n132), .C(\Queue[3][0] ), .D(n131), 
        .Z(n100) );
  OAI21M1P U248 ( .A(n143), .B(n134), .C(n100), .Z(n476) );
  AOI22M1P U249 ( .A(\Queue[2][1] ), .B(n132), .C(n131), .D(\Queue[3][1] ), 
        .Z(n101) );
  OAI21M1P U250 ( .A(n145), .B(n134), .C(n101), .Z(n477) );
  AOI22M1P U251 ( .A(\Queue[2][2] ), .B(n132), .C(n131), .D(\Queue[3][2] ), 
        .Z(n102) );
  OAI21M1P U252 ( .A(n147), .B(n134), .C(n102), .Z(n478) );
  AOI22M1P U253 ( .A(\Queue[2][3] ), .B(n132), .C(n131), .D(\Queue[3][3] ), 
        .Z(n103) );
  OAI21M1P U254 ( .A(n149), .B(n134), .C(n103), .Z(n479) );
  AOI22M1P U255 ( .A(\Queue[2][4] ), .B(n132), .C(n131), .D(\Queue[3][4] ), 
        .Z(n104) );
  OAI21M1P U256 ( .A(n151), .B(n134), .C(n104), .Z(n480) );
  AOI22M1P U257 ( .A(\Queue[2][5] ), .B(n132), .C(n131), .D(\Queue[3][5] ), 
        .Z(n105) );
  OAI21M1P U258 ( .A(n153), .B(n134), .C(n105), .Z(n481) );
  AOI22M1P U259 ( .A(\Queue[2][6] ), .B(n132), .C(n131), .D(\Queue[3][6] ), 
        .Z(n106) );
  OAI21M1P U260 ( .A(n155), .B(n134), .C(n106), .Z(n482) );
  AOI22M1P U261 ( .A(\Queue[2][7] ), .B(n132), .C(n131), .D(\Queue[3][7] ), 
        .Z(n107) );
  OAI21M1P U262 ( .A(n157), .B(n134), .C(n107), .Z(n483) );
  AOI22M1P U263 ( .A(\Queue[2][8] ), .B(n132), .C(n131), .D(\Queue[3][8] ), 
        .Z(n108) );
  OAI21M1P U264 ( .A(n159), .B(n134), .C(n108), .Z(n484) );
  AOI22M1P U265 ( .A(\Queue[2][9] ), .B(n132), .C(n131), .D(\Queue[3][9] ), 
        .Z(n109) );
  OAI21M1P U266 ( .A(n161), .B(n134), .C(n109), .Z(n485) );
  AOI22M1P U267 ( .A(\Queue[2][10] ), .B(n132), .C(n131), .D(\Queue[3][10] ), 
        .Z(n110) );
  OAI21M1P U268 ( .A(n163), .B(n134), .C(n110), .Z(n486) );
  AOI22M1P U269 ( .A(\Queue[2][11] ), .B(n132), .C(n131), .D(\Queue[3][11] ), 
        .Z(n111) );
  OAI21M1P U270 ( .A(n165), .B(n134), .C(n111), .Z(n487) );
  AOI22M1P U271 ( .A(\Queue[2][12] ), .B(n132), .C(n131), .D(\Queue[3][12] ), 
        .Z(n112) );
  OAI21M1P U272 ( .A(n167), .B(n134), .C(n112), .Z(n488) );
  AOI22M1P U273 ( .A(\Queue[2][13] ), .B(n132), .C(n131), .D(\Queue[3][13] ), 
        .Z(n113) );
  OAI21M1P U274 ( .A(n169), .B(n134), .C(n113), .Z(n489) );
  AOI22M1P U275 ( .A(\Queue[2][14] ), .B(n132), .C(n131), .D(\Queue[3][14] ), 
        .Z(n114) );
  OAI21M1P U276 ( .A(n171), .B(n134), .C(n114), .Z(n490) );
  AOI22M1P U277 ( .A(\Queue[2][15] ), .B(n132), .C(n131), .D(\Queue[3][15] ), 
        .Z(n115) );
  OAI21M1P U278 ( .A(n173), .B(n134), .C(n115), .Z(n491) );
  AOI22M1P U279 ( .A(\Queue[2][16] ), .B(n132), .C(n131), .D(\Queue[3][16] ), 
        .Z(n116) );
  OAI21M1P U280 ( .A(n175), .B(n134), .C(n116), .Z(n492) );
  AOI22M1P U281 ( .A(\Queue[2][17] ), .B(n132), .C(n131), .D(\Queue[3][17] ), 
        .Z(n117) );
  OAI21M1P U282 ( .A(n177), .B(n134), .C(n117), .Z(n493) );
  AOI22M1P U283 ( .A(\Queue[2][18] ), .B(n132), .C(n131), .D(\Queue[3][18] ), 
        .Z(n118) );
  OAI21M1P U284 ( .A(n179), .B(n134), .C(n118), .Z(n494) );
  AOI22M1P U285 ( .A(\Queue[2][19] ), .B(n132), .C(n131), .D(\Queue[3][19] ), 
        .Z(n119) );
  OAI21M1P U286 ( .A(n181), .B(n134), .C(n119), .Z(n495) );
  AOI22M1P U287 ( .A(\Queue[2][20] ), .B(n132), .C(n131), .D(\Queue[3][20] ), 
        .Z(n120) );
  OAI21M1P U288 ( .A(n183), .B(n134), .C(n120), .Z(n496) );
  AOI22M1P U289 ( .A(\Queue[2][21] ), .B(n132), .C(n131), .D(\Queue[3][21] ), 
        .Z(n121) );
  OAI21M1P U290 ( .A(n185), .B(n134), .C(n121), .Z(n497) );
  AOI22M1P U291 ( .A(\Queue[2][22] ), .B(n132), .C(n131), .D(\Queue[3][22] ), 
        .Z(n122) );
  OAI21M1P U292 ( .A(n187), .B(n134), .C(n122), .Z(n498) );
  AOI22M1P U293 ( .A(\Queue[2][23] ), .B(n132), .C(n131), .D(\Queue[3][23] ), 
        .Z(n123) );
  OAI21M1P U294 ( .A(n189), .B(n134), .C(n123), .Z(n499) );
  AOI22M1P U295 ( .A(\Queue[2][24] ), .B(n132), .C(n131), .D(\Queue[3][24] ), 
        .Z(n124) );
  OAI21M1P U296 ( .A(n191), .B(n134), .C(n124), .Z(n500) );
  AOI22M1P U297 ( .A(\Queue[2][25] ), .B(n132), .C(n131), .D(\Queue[3][25] ), 
        .Z(n125) );
  OAI21M1P U298 ( .A(n193), .B(n134), .C(n125), .Z(n501) );
  AOI22M1P U299 ( .A(\Queue[2][26] ), .B(n132), .C(n131), .D(\Queue[3][26] ), 
        .Z(n126) );
  OAI21M1P U300 ( .A(n195), .B(n134), .C(n126), .Z(n502) );
  AOI22M1P U301 ( .A(\Queue[2][27] ), .B(n132), .C(n131), .D(\Queue[3][27] ), 
        .Z(n127) );
  OAI21M1P U302 ( .A(n197), .B(n134), .C(n127), .Z(n503) );
  AOI22M1P U303 ( .A(\Queue[2][28] ), .B(n132), .C(n131), .D(\Queue[3][28] ), 
        .Z(n128) );
  OAI21M1P U304 ( .A(n199), .B(n134), .C(n128), .Z(n504) );
  AOI22M1P U305 ( .A(\Queue[2][29] ), .B(n132), .C(n131), .D(\Queue[3][29] ), 
        .Z(n129) );
  OAI21M1P U306 ( .A(n201), .B(n134), .C(n129), .Z(n505) );
  AOI22M1P U307 ( .A(\Queue[2][30] ), .B(n132), .C(n131), .D(\Queue[3][30] ), 
        .Z(n130) );
  OAI21M1P U308 ( .A(n203), .B(n134), .C(n130), .Z(n506) );
  AOI22M1P U309 ( .A(\Queue[2][31] ), .B(n132), .C(n131), .D(\Queue[3][31] ), 
        .Z(n133) );
  OAI21M1P U310 ( .A(n208), .B(n134), .C(n133), .Z(n507) );
  OA21M1P U311 ( .A(n138), .B(n139), .C(Rst_n), .Z(n135) );
  AOI22M1P U312 ( .A(\Queue[3][0] ), .B(n10), .C(n204), .D(\Queue[4][0] ), .Z(
        n142) );
  OAI21M1P U313 ( .A(n143), .B(n207), .C(n142), .Z(n508) );
  AOI22M1P U314 ( .A(\Queue[3][1] ), .B(n10), .C(n204), .D(\Queue[4][1] ), .Z(
        n144) );
  OAI21M1P U315 ( .A(n145), .B(n207), .C(n144), .Z(n509) );
  AOI22M1P U316 ( .A(\Queue[3][2] ), .B(n10), .C(n204), .D(\Queue[4][2] ), .Z(
        n146) );
  OAI21M1P U317 ( .A(n147), .B(n207), .C(n146), .Z(n510) );
  AOI22M1P U318 ( .A(\Queue[3][3] ), .B(n10), .C(n204), .D(\Queue[4][3] ), .Z(
        n148) );
  OAI21M1P U319 ( .A(n149), .B(n207), .C(n148), .Z(n511) );
  AOI22M1P U320 ( .A(\Queue[3][4] ), .B(n10), .C(n204), .D(\Queue[4][4] ), .Z(
        n150) );
  OAI21M1P U321 ( .A(n151), .B(n207), .C(n150), .Z(n512) );
  AOI22M1P U322 ( .A(\Queue[3][5] ), .B(n10), .C(n204), .D(\Queue[4][5] ), .Z(
        n152) );
  OAI21M1P U323 ( .A(n153), .B(n207), .C(n152), .Z(n513) );
  AOI22M1P U324 ( .A(\Queue[3][6] ), .B(n10), .C(n204), .D(\Queue[4][6] ), .Z(
        n154) );
  OAI21M1P U325 ( .A(n155), .B(n207), .C(n154), .Z(n514) );
  AOI22M1P U326 ( .A(\Queue[3][7] ), .B(n10), .C(n204), .D(\Queue[4][7] ), .Z(
        n156) );
  OAI21M1P U327 ( .A(n157), .B(n207), .C(n156), .Z(n515) );
  AOI22M1P U328 ( .A(\Queue[3][8] ), .B(n10), .C(n204), .D(\Queue[4][8] ), .Z(
        n158) );
  OAI21M1P U329 ( .A(n159), .B(n207), .C(n158), .Z(n516) );
  AOI22M1P U330 ( .A(\Queue[3][9] ), .B(n10), .C(n204), .D(\Queue[4][9] ), .Z(
        n160) );
  OAI21M1P U331 ( .A(n161), .B(n207), .C(n160), .Z(n517) );
  AOI22M1P U332 ( .A(\Queue[3][10] ), .B(n10), .C(n204), .D(\Queue[4][10] ), 
        .Z(n162) );
  OAI21M1P U333 ( .A(n163), .B(n207), .C(n162), .Z(n518) );
  AOI22M1P U334 ( .A(\Queue[3][11] ), .B(n10), .C(n204), .D(\Queue[4][11] ), 
        .Z(n164) );
  OAI21M1P U335 ( .A(n165), .B(n207), .C(n164), .Z(n519) );
  AOI22M1P U336 ( .A(\Queue[3][12] ), .B(n10), .C(n204), .D(\Queue[4][12] ), 
        .Z(n166) );
  OAI21M1P U337 ( .A(n167), .B(n207), .C(n166), .Z(n520) );
  AOI22M1P U338 ( .A(\Queue[3][13] ), .B(n10), .C(n204), .D(\Queue[4][13] ), 
        .Z(n168) );
  OAI21M1P U339 ( .A(n169), .B(n207), .C(n168), .Z(n521) );
  AOI22M1P U340 ( .A(\Queue[3][14] ), .B(n10), .C(n204), .D(\Queue[4][14] ), 
        .Z(n170) );
  OAI21M1P U341 ( .A(n171), .B(n207), .C(n170), .Z(n522) );
  AOI22M1P U342 ( .A(\Queue[3][15] ), .B(n10), .C(n204), .D(\Queue[4][15] ), 
        .Z(n172) );
  OAI21M1P U343 ( .A(n173), .B(n207), .C(n172), .Z(n523) );
  AOI22M1P U344 ( .A(\Queue[3][16] ), .B(n10), .C(n204), .D(\Queue[4][16] ), 
        .Z(n174) );
  OAI21M1P U345 ( .A(n175), .B(n207), .C(n174), .Z(n524) );
  AOI22M1P U346 ( .A(\Queue[3][17] ), .B(n10), .C(n204), .D(\Queue[4][17] ), 
        .Z(n176) );
  OAI21M1P U347 ( .A(n177), .B(n207), .C(n176), .Z(n525) );
  AOI22M1P U348 ( .A(\Queue[3][18] ), .B(n10), .C(n204), .D(\Queue[4][18] ), 
        .Z(n178) );
  OAI21M1P U349 ( .A(n179), .B(n207), .C(n178), .Z(n526) );
  AOI22M1P U350 ( .A(\Queue[3][19] ), .B(n10), .C(n204), .D(\Queue[4][19] ), 
        .Z(n180) );
  OAI21M1P U351 ( .A(n181), .B(n207), .C(n180), .Z(n527) );
  AOI22M1P U352 ( .A(\Queue[3][20] ), .B(n11), .C(n204), .D(\Queue[4][20] ), 
        .Z(n182) );
  OAI21M1P U353 ( .A(n183), .B(n207), .C(n182), .Z(n528) );
  AOI22M1P U354 ( .A(\Queue[3][21] ), .B(n11), .C(n204), .D(\Queue[4][21] ), 
        .Z(n184) );
  OAI21M1P U355 ( .A(n185), .B(n207), .C(n184), .Z(n529) );
  AOI22M1P U356 ( .A(\Queue[3][22] ), .B(n11), .C(n204), .D(\Queue[4][22] ), 
        .Z(n186) );
  OAI21M1P U357 ( .A(n187), .B(n207), .C(n186), .Z(n530) );
  AOI22M1P U358 ( .A(\Queue[3][23] ), .B(n11), .C(n204), .D(\Queue[4][23] ), 
        .Z(n188) );
  OAI21M1P U359 ( .A(n189), .B(n207), .C(n188), .Z(n531) );
  AOI22M1P U360 ( .A(\Queue[3][24] ), .B(n11), .C(n204), .D(\Queue[4][24] ), 
        .Z(n190) );
  OAI21M1P U361 ( .A(n191), .B(n207), .C(n190), .Z(n532) );
  AOI22M1P U362 ( .A(\Queue[3][25] ), .B(n11), .C(n204), .D(\Queue[4][25] ), 
        .Z(n192) );
  OAI21M1P U363 ( .A(n193), .B(n207), .C(n192), .Z(n533) );
  AOI22M1P U364 ( .A(\Queue[3][26] ), .B(n11), .C(n204), .D(\Queue[4][26] ), 
        .Z(n194) );
  OAI21M1P U365 ( .A(n195), .B(n207), .C(n194), .Z(n534) );
  AOI22M1P U366 ( .A(\Queue[3][27] ), .B(n11), .C(n204), .D(\Queue[4][27] ), 
        .Z(n196) );
  OAI21M1P U367 ( .A(n197), .B(n207), .C(n196), .Z(n535) );
  AOI22M1P U368 ( .A(\Queue[3][28] ), .B(n11), .C(n204), .D(\Queue[4][28] ), 
        .Z(n198) );
  OAI21M1P U369 ( .A(n199), .B(n207), .C(n198), .Z(n536) );
  AOI22M1P U370 ( .A(\Queue[3][29] ), .B(n11), .C(n204), .D(\Queue[4][29] ), 
        .Z(n200) );
  OAI21M1P U371 ( .A(n201), .B(n207), .C(n200), .Z(n537) );
  AOI22M1P U372 ( .A(\Queue[3][30] ), .B(n10), .C(n204), .D(\Queue[4][30] ), 
        .Z(n202) );
  OAI21M1P U373 ( .A(n203), .B(n207), .C(n202), .Z(n538) );
  AOI22M1P U374 ( .A(\Queue[3][31] ), .B(n11), .C(n204), .D(\Queue[4][31] ), 
        .Z(n206) );
  OAI21M1P U375 ( .A(n208), .B(n207), .C(n206), .Z(n539) );
  N1M1P U376 ( .A(n540), .Z(Empty) );
  AOI22M1P U377 ( .A(n375), .B(n374), .C(n373), .D(Empty), .Z(n541) );
endmodule


module Packet_Queue_6 ( Clk_r, Rst_n, Packet_In, Read_Ack, Write_Ack, 
        Packet_Out, Empty, Full );
  input [31:0] Packet_In;
  output [31:0] Packet_Out;
  input Clk_r, Rst_n, Read_Ack, Write_Ack;
  output Empty, Full;
  wire   \Queue[4][31] , \Queue[4][30] , \Queue[4][29] , \Queue[4][28] ,
         \Queue[4][27] , \Queue[4][26] , \Queue[4][25] , \Queue[4][24] ,
         \Queue[4][23] , \Queue[4][22] , \Queue[4][21] , \Queue[4][20] ,
         \Queue[4][19] , \Queue[4][18] , \Queue[4][17] , \Queue[4][16] ,
         \Queue[4][15] , \Queue[4][14] , \Queue[4][13] , \Queue[4][12] ,
         \Queue[4][11] , \Queue[4][10] , \Queue[4][9] , \Queue[4][8] ,
         \Queue[4][7] , \Queue[4][6] , \Queue[4][5] , \Queue[4][4] ,
         \Queue[4][3] , \Queue[4][2] , \Queue[4][1] , \Queue[4][0] ,
         \Queue[3][31] , \Queue[3][30] , \Queue[3][29] , \Queue[3][28] ,
         \Queue[3][27] , \Queue[3][26] , \Queue[3][25] , \Queue[3][24] ,
         \Queue[3][23] , \Queue[3][22] , \Queue[3][21] , \Queue[3][20] ,
         \Queue[3][19] , \Queue[3][18] , \Queue[3][17] , \Queue[3][16] ,
         \Queue[3][15] , \Queue[3][14] , \Queue[3][13] , \Queue[3][12] ,
         \Queue[3][11] , \Queue[3][10] , \Queue[3][9] , \Queue[3][8] ,
         \Queue[3][7] , \Queue[3][6] , \Queue[3][5] , \Queue[3][4] ,
         \Queue[3][3] , \Queue[3][2] , \Queue[3][1] , \Queue[3][0] ,
         \Queue[2][31] , \Queue[2][30] , \Queue[2][29] , \Queue[2][28] ,
         \Queue[2][27] , \Queue[2][26] , \Queue[2][25] , \Queue[2][24] ,
         \Queue[2][23] , \Queue[2][22] , \Queue[2][21] , \Queue[2][20] ,
         \Queue[2][19] , \Queue[2][18] , \Queue[2][17] , \Queue[2][16] ,
         \Queue[2][15] , \Queue[2][14] , \Queue[2][13] , \Queue[2][12] ,
         \Queue[2][11] , \Queue[2][10] , \Queue[2][9] , \Queue[2][8] ,
         \Queue[2][7] , \Queue[2][6] , \Queue[2][5] , \Queue[2][4] ,
         \Queue[2][3] , \Queue[2][2] , \Queue[2][1] , \Queue[2][0] ,
         \Queue[1][31] , \Queue[1][30] , \Queue[1][29] , \Queue[1][28] ,
         \Queue[1][27] , \Queue[1][26] , \Queue[1][25] , \Queue[1][24] ,
         \Queue[1][23] , \Queue[1][22] , \Queue[1][21] , \Queue[1][20] ,
         \Queue[1][19] , \Queue[1][18] , \Queue[1][17] , \Queue[1][16] ,
         \Queue[1][15] , \Queue[1][14] , \Queue[1][13] , \Queue[1][12] ,
         \Queue[1][11] , \Queue[1][10] , \Queue[1][9] , \Queue[1][8] ,
         \Queue[1][7] , \Queue[1][6] , \Queue[1][5] , \Queue[1][4] ,
         \Queue[1][3] , \Queue[1][2] , \Queue[1][1] , \Queue[1][0] , n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547;
  wire   [2:0] Count;

  FDN2QM1P \Count_reg[0]  ( .D(n382), .CPN(Clk_r), .CD(Rst_n), .Q(Count[0]) );
  FDN2QM1P \Count_reg[1]  ( .D(n383), .CPN(Clk_r), .CD(Rst_n), .Q(Count[1]) );
  FDN2QM1P \Count_reg[2]  ( .D(n384), .CPN(Clk_r), .CD(Rst_n), .Q(Count[2]) );
  FDN1QM1P \Queue_reg[4][30]  ( .D(n416), .CPN(Clk_r), .Q(\Queue[4][30] ) );
  FDN1QM1P \Queue_reg[3][30]  ( .D(n544), .CPN(Clk_r), .Q(\Queue[3][30] ) );
  FDN1QM1P \Queue_reg[2][30]  ( .D(n512), .CPN(Clk_r), .Q(\Queue[2][30] ) );
  FDN1QM1P \Queue_reg[4][29]  ( .D(n415), .CPN(Clk_r), .Q(\Queue[4][29] ) );
  FDN1QM1P \Queue_reg[3][29]  ( .D(n543), .CPN(Clk_r), .Q(\Queue[3][29] ) );
  FDN1QM1P \Queue_reg[2][29]  ( .D(n511), .CPN(Clk_r), .Q(\Queue[2][29] ) );
  FDN1QM1P \Queue_reg[4][28]  ( .D(n414), .CPN(Clk_r), .Q(\Queue[4][28] ) );
  FDN1QM1P \Queue_reg[3][28]  ( .D(n542), .CPN(Clk_r), .Q(\Queue[3][28] ) );
  FDN1QM1P \Queue_reg[2][28]  ( .D(n510), .CPN(Clk_r), .Q(\Queue[2][28] ) );
  FDN1QM1P \Queue_reg[4][27]  ( .D(n413), .CPN(Clk_r), .Q(\Queue[4][27] ) );
  FDN1QM1P \Queue_reg[3][27]  ( .D(n541), .CPN(Clk_r), .Q(\Queue[3][27] ) );
  FDN1QM1P \Queue_reg[2][27]  ( .D(n509), .CPN(Clk_r), .Q(\Queue[2][27] ) );
  FDN1QM1P \Queue_reg[4][26]  ( .D(n412), .CPN(Clk_r), .Q(\Queue[4][26] ) );
  FDN1QM1P \Queue_reg[3][26]  ( .D(n540), .CPN(Clk_r), .Q(\Queue[3][26] ) );
  FDN1QM1P \Queue_reg[2][26]  ( .D(n508), .CPN(Clk_r), .Q(\Queue[2][26] ) );
  FDN1QM1P \Queue_reg[4][25]  ( .D(n411), .CPN(Clk_r), .Q(\Queue[4][25] ) );
  FDN1QM1P \Queue_reg[3][25]  ( .D(n539), .CPN(Clk_r), .Q(\Queue[3][25] ) );
  FDN1QM1P \Queue_reg[2][25]  ( .D(n507), .CPN(Clk_r), .Q(\Queue[2][25] ) );
  FDN1QM1P \Queue_reg[4][24]  ( .D(n410), .CPN(Clk_r), .Q(\Queue[4][24] ) );
  FDN1QM1P \Queue_reg[3][24]  ( .D(n538), .CPN(Clk_r), .Q(\Queue[3][24] ) );
  FDN1QM1P \Queue_reg[2][24]  ( .D(n506), .CPN(Clk_r), .Q(\Queue[2][24] ) );
  FDN1QM1P \Queue_reg[4][23]  ( .D(n409), .CPN(Clk_r), .Q(\Queue[4][23] ) );
  FDN1QM1P \Queue_reg[3][23]  ( .D(n537), .CPN(Clk_r), .Q(\Queue[3][23] ) );
  FDN1QM1P \Queue_reg[2][23]  ( .D(n505), .CPN(Clk_r), .Q(\Queue[2][23] ) );
  FDN1QM1P \Queue_reg[4][22]  ( .D(n408), .CPN(Clk_r), .Q(\Queue[4][22] ) );
  FDN1QM1P \Queue_reg[3][22]  ( .D(n536), .CPN(Clk_r), .Q(\Queue[3][22] ) );
  FDN1QM1P \Queue_reg[2][22]  ( .D(n504), .CPN(Clk_r), .Q(\Queue[2][22] ) );
  FDN1QM1P \Queue_reg[4][21]  ( .D(n407), .CPN(Clk_r), .Q(\Queue[4][21] ) );
  FDN1QM1P \Queue_reg[3][21]  ( .D(n535), .CPN(Clk_r), .Q(\Queue[3][21] ) );
  FDN1QM1P \Queue_reg[2][21]  ( .D(n503), .CPN(Clk_r), .Q(\Queue[2][21] ) );
  FDN1QM1P \Queue_reg[4][20]  ( .D(n406), .CPN(Clk_r), .Q(\Queue[4][20] ) );
  FDN1QM1P \Queue_reg[3][20]  ( .D(n534), .CPN(Clk_r), .Q(\Queue[3][20] ) );
  FDN1QM1P \Queue_reg[2][20]  ( .D(n502), .CPN(Clk_r), .Q(\Queue[2][20] ) );
  FDN1QM1P \Queue_reg[4][19]  ( .D(n405), .CPN(Clk_r), .Q(\Queue[4][19] ) );
  FDN1QM1P \Queue_reg[3][19]  ( .D(n533), .CPN(Clk_r), .Q(\Queue[3][19] ) );
  FDN1QM1P \Queue_reg[2][19]  ( .D(n501), .CPN(Clk_r), .Q(\Queue[2][19] ) );
  FDN1QM1P \Queue_reg[4][18]  ( .D(n404), .CPN(Clk_r), .Q(\Queue[4][18] ) );
  FDN1QM1P \Queue_reg[3][18]  ( .D(n532), .CPN(Clk_r), .Q(\Queue[3][18] ) );
  FDN1QM1P \Queue_reg[2][18]  ( .D(n500), .CPN(Clk_r), .Q(\Queue[2][18] ) );
  FDN1QM1P \Queue_reg[4][17]  ( .D(n403), .CPN(Clk_r), .Q(\Queue[4][17] ) );
  FDN1QM1P \Queue_reg[3][17]  ( .D(n531), .CPN(Clk_r), .Q(\Queue[3][17] ) );
  FDN1QM1P \Queue_reg[2][17]  ( .D(n499), .CPN(Clk_r), .Q(\Queue[2][17] ) );
  FDN1QM1P \Queue_reg[4][16]  ( .D(n402), .CPN(Clk_r), .Q(\Queue[4][16] ) );
  FDN1QM1P \Queue_reg[3][16]  ( .D(n530), .CPN(Clk_r), .Q(\Queue[3][16] ) );
  FDN1QM1P \Queue_reg[2][16]  ( .D(n498), .CPN(Clk_r), .Q(\Queue[2][16] ) );
  FDN1QM1P \Queue_reg[4][15]  ( .D(n401), .CPN(Clk_r), .Q(\Queue[4][15] ) );
  FDN1QM1P \Queue_reg[3][15]  ( .D(n529), .CPN(Clk_r), .Q(\Queue[3][15] ) );
  FDN1QM1P \Queue_reg[2][15]  ( .D(n497), .CPN(Clk_r), .Q(\Queue[2][15] ) );
  FDN1QM1P \Queue_reg[4][14]  ( .D(n400), .CPN(Clk_r), .Q(\Queue[4][14] ) );
  FDN1QM1P \Queue_reg[3][14]  ( .D(n528), .CPN(Clk_r), .Q(\Queue[3][14] ) );
  FDN1QM1P \Queue_reg[2][14]  ( .D(n496), .CPN(Clk_r), .Q(\Queue[2][14] ) );
  FDN1QM1P \Queue_reg[4][13]  ( .D(n399), .CPN(Clk_r), .Q(\Queue[4][13] ) );
  FDN1QM1P \Queue_reg[3][13]  ( .D(n527), .CPN(Clk_r), .Q(\Queue[3][13] ) );
  FDN1QM1P \Queue_reg[2][13]  ( .D(n495), .CPN(Clk_r), .Q(\Queue[2][13] ) );
  FDN1QM1P \Queue_reg[4][12]  ( .D(n398), .CPN(Clk_r), .Q(\Queue[4][12] ) );
  FDN1QM1P \Queue_reg[3][12]  ( .D(n526), .CPN(Clk_r), .Q(\Queue[3][12] ) );
  FDN1QM1P \Queue_reg[2][12]  ( .D(n494), .CPN(Clk_r), .Q(\Queue[2][12] ) );
  FDN1QM1P \Queue_reg[4][11]  ( .D(n397), .CPN(Clk_r), .Q(\Queue[4][11] ) );
  FDN1QM1P \Queue_reg[3][11]  ( .D(n525), .CPN(Clk_r), .Q(\Queue[3][11] ) );
  FDN1QM1P \Queue_reg[2][11]  ( .D(n493), .CPN(Clk_r), .Q(\Queue[2][11] ) );
  FDN1QM1P \Queue_reg[4][10]  ( .D(n396), .CPN(Clk_r), .Q(\Queue[4][10] ) );
  FDN1QM1P \Queue_reg[3][10]  ( .D(n524), .CPN(Clk_r), .Q(\Queue[3][10] ) );
  FDN1QM1P \Queue_reg[2][10]  ( .D(n492), .CPN(Clk_r), .Q(\Queue[2][10] ) );
  FDN1QM1P \Queue_reg[4][9]  ( .D(n395), .CPN(Clk_r), .Q(\Queue[4][9] ) );
  FDN1QM1P \Queue_reg[3][9]  ( .D(n523), .CPN(Clk_r), .Q(\Queue[3][9] ) );
  FDN1QM1P \Queue_reg[2][9]  ( .D(n491), .CPN(Clk_r), .Q(\Queue[2][9] ) );
  FDN1QM1P \Queue_reg[4][8]  ( .D(n394), .CPN(Clk_r), .Q(\Queue[4][8] ) );
  FDN1QM1P \Queue_reg[3][8]  ( .D(n522), .CPN(Clk_r), .Q(\Queue[3][8] ) );
  FDN1QM1P \Queue_reg[2][8]  ( .D(n490), .CPN(Clk_r), .Q(\Queue[2][8] ) );
  FDN1QM1P \Queue_reg[4][7]  ( .D(n393), .CPN(Clk_r), .Q(\Queue[4][7] ) );
  FDN1QM1P \Queue_reg[3][7]  ( .D(n521), .CPN(Clk_r), .Q(\Queue[3][7] ) );
  FDN1QM1P \Queue_reg[2][7]  ( .D(n489), .CPN(Clk_r), .Q(\Queue[2][7] ) );
  FDN1QM1P \Queue_reg[4][6]  ( .D(n392), .CPN(Clk_r), .Q(\Queue[4][6] ) );
  FDN1QM1P \Queue_reg[3][6]  ( .D(n520), .CPN(Clk_r), .Q(\Queue[3][6] ) );
  FDN1QM1P \Queue_reg[2][6]  ( .D(n488), .CPN(Clk_r), .Q(\Queue[2][6] ) );
  FDN1QM1P \Queue_reg[4][5]  ( .D(n391), .CPN(Clk_r), .Q(\Queue[4][5] ) );
  FDN1QM1P \Queue_reg[3][5]  ( .D(n519), .CPN(Clk_r), .Q(\Queue[3][5] ) );
  FDN1QM1P \Queue_reg[2][5]  ( .D(n487), .CPN(Clk_r), .Q(\Queue[2][5] ) );
  FDN1QM1P \Queue_reg[4][4]  ( .D(n390), .CPN(Clk_r), .Q(\Queue[4][4] ) );
  FDN1QM1P \Queue_reg[3][4]  ( .D(n518), .CPN(Clk_r), .Q(\Queue[3][4] ) );
  FDN1QM1P \Queue_reg[2][4]  ( .D(n486), .CPN(Clk_r), .Q(\Queue[2][4] ) );
  FDN1QM1P \Queue_reg[4][3]  ( .D(n389), .CPN(Clk_r), .Q(\Queue[4][3] ) );
  FDN1QM1P \Queue_reg[3][3]  ( .D(n517), .CPN(Clk_r), .Q(\Queue[3][3] ) );
  FDN1QM1P \Queue_reg[2][3]  ( .D(n485), .CPN(Clk_r), .Q(\Queue[2][3] ) );
  FDN1QM1P \Queue_reg[4][2]  ( .D(n388), .CPN(Clk_r), .Q(\Queue[4][2] ) );
  FDN1QM1P \Queue_reg[3][2]  ( .D(n516), .CPN(Clk_r), .Q(\Queue[3][2] ) );
  FDN1QM1P \Queue_reg[2][2]  ( .D(n484), .CPN(Clk_r), .Q(\Queue[2][2] ) );
  FDN1QM1P \Queue_reg[4][1]  ( .D(n387), .CPN(Clk_r), .Q(\Queue[4][1] ) );
  FDN1QM1P \Queue_reg[3][1]  ( .D(n515), .CPN(Clk_r), .Q(\Queue[3][1] ) );
  FDN1QM1P \Queue_reg[2][1]  ( .D(n483), .CPN(Clk_r), .Q(\Queue[2][1] ) );
  FDN1QM1P \Queue_reg[4][0]  ( .D(n386), .CPN(Clk_r), .Q(\Queue[4][0] ) );
  FDN1QM1P \Queue_reg[3][0]  ( .D(n514), .CPN(Clk_r), .Q(\Queue[3][0] ) );
  FDN1QM1P \Queue_reg[2][0]  ( .D(n482), .CPN(Clk_r), .Q(\Queue[2][0] ) );
  FDN1QM1P \Queue_reg[4][31]  ( .D(n385), .CPN(Clk_r), .Q(\Queue[4][31] ) );
  FDN1QM1P \Queue_reg[3][31]  ( .D(n545), .CPN(Clk_r), .Q(\Queue[3][31] ) );
  FDN1QM1P \Queue_reg[2][31]  ( .D(n513), .CPN(Clk_r), .Q(\Queue[2][31] ) );
  FDN2QM1P Full_reg ( .D(n417), .CPN(Clk_r), .CD(Rst_n), .Q(Full) );
  FDN1QM1P \Queue_reg[1][31]  ( .D(n449), .CPN(Clk_r), .Q(\Queue[1][31] ) );
  FDN1QM1P \Queue_reg[0][31]  ( .D(n481), .CPN(Clk_r), .Q(Packet_Out[31]) );
  FDN1QM1P \Queue_reg[1][30]  ( .D(n448), .CPN(Clk_r), .Q(\Queue[1][30] ) );
  FDN1QM1P \Queue_reg[0][30]  ( .D(n480), .CPN(Clk_r), .Q(Packet_Out[30]) );
  FDN1QM1P \Queue_reg[1][29]  ( .D(n447), .CPN(Clk_r), .Q(\Queue[1][29] ) );
  FDN1QM1P \Queue_reg[0][29]  ( .D(n479), .CPN(Clk_r), .Q(Packet_Out[29]) );
  FDN1QM1P \Queue_reg[1][28]  ( .D(n446), .CPN(Clk_r), .Q(\Queue[1][28] ) );
  FDN1QM1P \Queue_reg[0][28]  ( .D(n478), .CPN(Clk_r), .Q(Packet_Out[28]) );
  FDN1QM1P \Queue_reg[1][27]  ( .D(n445), .CPN(Clk_r), .Q(\Queue[1][27] ) );
  FDN1QM1P \Queue_reg[0][27]  ( .D(n477), .CPN(Clk_r), .Q(Packet_Out[27]) );
  FDN1QM1P \Queue_reg[1][26]  ( .D(n444), .CPN(Clk_r), .Q(\Queue[1][26] ) );
  FDN1QM1P \Queue_reg[0][26]  ( .D(n476), .CPN(Clk_r), .Q(Packet_Out[26]) );
  FDN1QM1P \Queue_reg[1][25]  ( .D(n443), .CPN(Clk_r), .Q(\Queue[1][25] ) );
  FDN1QM1P \Queue_reg[0][25]  ( .D(n475), .CPN(Clk_r), .Q(Packet_Out[25]) );
  FDN1QM1P \Queue_reg[1][24]  ( .D(n442), .CPN(Clk_r), .Q(\Queue[1][24] ) );
  FDN1QM1P \Queue_reg[0][24]  ( .D(n474), .CPN(Clk_r), .Q(Packet_Out[24]) );
  FDN1QM1P \Queue_reg[1][23]  ( .D(n441), .CPN(Clk_r), .Q(\Queue[1][23] ) );
  FDN1QM1P \Queue_reg[0][23]  ( .D(n473), .CPN(Clk_r), .Q(Packet_Out[23]) );
  FDN1QM1P \Queue_reg[1][22]  ( .D(n440), .CPN(Clk_r), .Q(\Queue[1][22] ) );
  FDN1QM1P \Queue_reg[0][22]  ( .D(n472), .CPN(Clk_r), .Q(Packet_Out[22]) );
  FDN1QM1P \Queue_reg[1][21]  ( .D(n439), .CPN(Clk_r), .Q(\Queue[1][21] ) );
  FDN1QM1P \Queue_reg[0][21]  ( .D(n471), .CPN(Clk_r), .Q(Packet_Out[21]) );
  FDN1QM1P \Queue_reg[1][20]  ( .D(n438), .CPN(Clk_r), .Q(\Queue[1][20] ) );
  FDN1QM1P \Queue_reg[0][20]  ( .D(n470), .CPN(Clk_r), .Q(Packet_Out[20]) );
  FDN1QM1P \Queue_reg[1][19]  ( .D(n437), .CPN(Clk_r), .Q(\Queue[1][19] ) );
  FDN1QM1P \Queue_reg[0][19]  ( .D(n469), .CPN(Clk_r), .Q(Packet_Out[19]) );
  FDN1QM1P \Queue_reg[1][18]  ( .D(n436), .CPN(Clk_r), .Q(\Queue[1][18] ) );
  FDN1QM1P \Queue_reg[0][18]  ( .D(n468), .CPN(Clk_r), .Q(Packet_Out[18]) );
  FDN1QM1P \Queue_reg[1][17]  ( .D(n435), .CPN(Clk_r), .Q(\Queue[1][17] ) );
  FDN1QM1P \Queue_reg[0][17]  ( .D(n467), .CPN(Clk_r), .Q(Packet_Out[17]) );
  FDN1QM1P \Queue_reg[1][16]  ( .D(n434), .CPN(Clk_r), .Q(\Queue[1][16] ) );
  FDN1QM1P \Queue_reg[0][16]  ( .D(n466), .CPN(Clk_r), .Q(Packet_Out[16]) );
  FDN1QM1P \Queue_reg[1][15]  ( .D(n433), .CPN(Clk_r), .Q(\Queue[1][15] ) );
  FDN1QM1P \Queue_reg[0][15]  ( .D(n465), .CPN(Clk_r), .Q(Packet_Out[15]) );
  FDN1QM1P \Queue_reg[1][14]  ( .D(n432), .CPN(Clk_r), .Q(\Queue[1][14] ) );
  FDN1QM1P \Queue_reg[0][14]  ( .D(n464), .CPN(Clk_r), .Q(Packet_Out[14]) );
  FDN1QM1P \Queue_reg[1][13]  ( .D(n431), .CPN(Clk_r), .Q(\Queue[1][13] ) );
  FDN1QM1P \Queue_reg[0][13]  ( .D(n463), .CPN(Clk_r), .Q(Packet_Out[13]) );
  FDN1QM1P \Queue_reg[1][12]  ( .D(n430), .CPN(Clk_r), .Q(\Queue[1][12] ) );
  FDN1QM1P \Queue_reg[0][12]  ( .D(n462), .CPN(Clk_r), .Q(Packet_Out[12]) );
  FDN1QM1P \Queue_reg[1][11]  ( .D(n429), .CPN(Clk_r), .Q(\Queue[1][11] ) );
  FDN1QM1P \Queue_reg[0][11]  ( .D(n461), .CPN(Clk_r), .Q(Packet_Out[11]) );
  FDN1QM1P \Queue_reg[1][10]  ( .D(n428), .CPN(Clk_r), .Q(\Queue[1][10] ) );
  FDN1QM1P \Queue_reg[0][10]  ( .D(n460), .CPN(Clk_r), .Q(Packet_Out[10]) );
  FDN1QM1P \Queue_reg[1][9]  ( .D(n427), .CPN(Clk_r), .Q(\Queue[1][9] ) );
  FDN1QM1P \Queue_reg[0][9]  ( .D(n459), .CPN(Clk_r), .Q(Packet_Out[9]) );
  FDN1QM1P \Queue_reg[1][8]  ( .D(n426), .CPN(Clk_r), .Q(\Queue[1][8] ) );
  FDN1QM1P \Queue_reg[0][8]  ( .D(n458), .CPN(Clk_r), .Q(Packet_Out[8]) );
  FDN1QM1P \Queue_reg[1][7]  ( .D(n425), .CPN(Clk_r), .Q(\Queue[1][7] ) );
  FDN1QM1P \Queue_reg[0][7]  ( .D(n457), .CPN(Clk_r), .Q(Packet_Out[7]) );
  FDN1QM1P \Queue_reg[1][6]  ( .D(n424), .CPN(Clk_r), .Q(\Queue[1][6] ) );
  FDN1QM1P \Queue_reg[0][6]  ( .D(n456), .CPN(Clk_r), .Q(Packet_Out[6]) );
  FDN1QM1P \Queue_reg[1][5]  ( .D(n423), .CPN(Clk_r), .Q(\Queue[1][5] ) );
  FDN1QM1P \Queue_reg[0][5]  ( .D(n455), .CPN(Clk_r), .Q(Packet_Out[5]) );
  FDN1QM1P \Queue_reg[1][4]  ( .D(n422), .CPN(Clk_r), .Q(\Queue[1][4] ) );
  FDN1QM1P \Queue_reg[0][4]  ( .D(n454), .CPN(Clk_r), .Q(Packet_Out[4]) );
  FDN1QM1P \Queue_reg[1][3]  ( .D(n421), .CPN(Clk_r), .Q(\Queue[1][3] ) );
  FDN1QM1P \Queue_reg[0][3]  ( .D(n453), .CPN(Clk_r), .Q(Packet_Out[3]) );
  FDN1QM1P \Queue_reg[1][2]  ( .D(n420), .CPN(Clk_r), .Q(\Queue[1][2] ) );
  FDN1QM1P \Queue_reg[0][2]  ( .D(n452), .CPN(Clk_r), .Q(Packet_Out[2]) );
  FDN1QM1P \Queue_reg[1][1]  ( .D(n419), .CPN(Clk_r), .Q(\Queue[1][1] ) );
  FDN1QM1P \Queue_reg[0][1]  ( .D(n451), .CPN(Clk_r), .Q(Packet_Out[1]) );
  FDN1QM1P \Queue_reg[1][0]  ( .D(n418), .CPN(Clk_r), .Q(\Queue[1][0] ) );
  FDN1QM1P \Queue_reg[0][0]  ( .D(n450), .CPN(Clk_r), .Q(Packet_Out[0]) );
  FDN2QM1P Empty_reg ( .D(n547), .CPN(Clk_r), .CD(Rst_n), .Q(n546) );
  BUFM2P U3 ( .A(n67), .Z(n43) );
  N1M2P U4 ( .A(n72), .Z(n104) );
  BUFM2P U5 ( .A(n67), .Z(n42) );
  BUFM1P U6 ( .A(n141), .Z(n49) );
  BUFM1P U7 ( .A(n375), .Z(n52) );
  BUFM2P U8 ( .A(n141), .Z(n48) );
  ND2M2P U9 ( .A(n7), .B(n8), .Z(n50) );
  BUFM2P U10 ( .A(n375), .Z(n51) );
  AOI21M8P U11 ( .A(n41), .B(n146), .C(n147), .Z(n140) );
  ND2M1P U12 ( .A(Read_Ack), .B(Rst_n), .Z(n147) );
  AOI21M3P U13 ( .A(n41), .B(n109), .C(n147), .Z(n68) );
  AOI21M3P U14 ( .A(n41), .B(n148), .C(n147), .Z(n374) );
  NR2FM3P U15 ( .A(n71), .B(n61), .Z(n60) );
  AOI21M3P U16 ( .A(n41), .B(n381), .C(n147), .Z(n105) );
  BUFM1P U17 ( .A(n107), .Z(n46) );
  N1M2P U18 ( .A(n41), .Z(n108) );
  NR3M1P U19 ( .A(Count[0]), .B(Count[1]), .C(n59), .Z(n148) );
  BUFM6P U20 ( .A(Write_Ack), .Z(n41) );
  ND2BNM2P U21 ( .B(n3), .A(n4), .Z(n377) );
  N1M2P U22 ( .A(n58), .Z(n145) );
  N1M1P U23 ( .A(n148), .Z(n61) );
  NR3M1P U24 ( .A(Count[2]), .B(n63), .C(n62), .Z(n146) );
  NR3M1P U25 ( .A(n63), .B(Count[2]), .C(Count[1]), .Z(n381) );
  NR3M1P U26 ( .A(Count[0]), .B(Count[2]), .C(n62), .Z(n109) );
  N1M1P U27 ( .A(Count[0]), .Z(n63) );
  N1M1P U28 ( .A(Count[1]), .Z(n62) );
  N1M1P U29 ( .A(Count[2]), .Z(n59) );
  BUFM2P U30 ( .A(n69), .Z(n45) );
  NR2FM2P U31 ( .A(Read_Ack), .B(n108), .Z(n58) );
  ND2M2P U32 ( .A(n58), .B(Rst_n), .Z(n71) );
  OAI21M2P U33 ( .A(n71), .B(n70), .C(n147), .Z(n72) );
  OAI211M1P U34 ( .A(n381), .B(n143), .C(n41), .D(n72), .Z(n107) );
  BUFM2P U35 ( .A(n69), .Z(n44) );
  N1M1P U36 ( .A(Read_Ack), .Z(n143) );
  N1M1P U37 ( .A(Packet_In[2]), .Z(n153) );
  N1M1P U38 ( .A(Packet_In[1]), .Z(n151) );
  N1M1P U39 ( .A(Packet_In[7]), .Z(n163) );
  N1M1P U40 ( .A(Packet_In[6]), .Z(n161) );
  N1M1P U41 ( .A(Packet_In[16]), .Z(n181) );
  N1M1P U42 ( .A(Packet_In[28]), .Z(n205) );
  N1M1P U43 ( .A(Packet_In[11]), .Z(n171) );
  N1M1P U44 ( .A(Packet_In[29]), .Z(n207) );
  N1M1P U45 ( .A(Packet_In[13]), .Z(n175) );
  N1M1P U46 ( .A(Packet_In[15]), .Z(n179) );
  N1M1P U47 ( .A(Packet_In[24]), .Z(n197) );
  N1M1P U48 ( .A(Packet_In[31]), .Z(n378) );
  N1M1P U49 ( .A(Packet_In[26]), .Z(n201) );
  N1M1P U50 ( .A(Packet_In[27]), .Z(n203) );
  N1M1P U51 ( .A(Packet_In[0]), .Z(n149) );
  N1M1P U52 ( .A(Packet_In[23]), .Z(n195) );
  N1M1P U53 ( .A(Packet_In[30]), .Z(n373) );
  N1M1P U54 ( .A(Packet_In[9]), .Z(n167) );
  N1M1P U55 ( .A(Packet_In[25]), .Z(n199) );
  N1M1P U56 ( .A(Packet_In[10]), .Z(n169) );
  N1M1P U57 ( .A(Packet_In[12]), .Z(n173) );
  N1M1P U58 ( .A(Packet_In[4]), .Z(n157) );
  N1M1P U59 ( .A(Packet_In[8]), .Z(n165) );
  N1M1P U60 ( .A(Packet_In[20]), .Z(n189) );
  N1M1P U61 ( .A(Packet_In[19]), .Z(n187) );
  N1M1P U62 ( .A(Packet_In[3]), .Z(n155) );
  N1M1P U63 ( .A(Packet_In[21]), .Z(n191) );
  N1M1P U64 ( .A(Packet_In[17]), .Z(n183) );
  N1M1P U65 ( .A(Packet_In[18]), .Z(n185) );
  N1M1P U66 ( .A(Packet_In[5]), .Z(n159) );
  N1M1P U67 ( .A(Packet_In[14]), .Z(n177) );
  N1M1P U68 ( .A(Packet_In[22]), .Z(n193) );
  BUFM2P U69 ( .A(n107), .Z(n47) );
  OA21M1P U70 ( .A(n145), .B(n381), .C(Rst_n), .Z(n64) );
  ND2BNM1P U71 ( .B(n146), .A(n5), .Z(n4) );
  OAI21M1P U72 ( .A(n149), .B(n45), .C(n65), .Z(n418) );
  AOI22M1P U73 ( .A(\Queue[2][0] ), .B(n68), .C(\Queue[1][0] ), .D(n42), .Z(
        n65) );
  AOI22M1P U74 ( .A(\Queue[2][1] ), .B(n48), .C(n140), .D(\Queue[3][1] ), .Z(
        n110) );
  N1M1P U75 ( .A(n145), .Z(n5) );
  OAI211M1P U76 ( .A(n148), .B(n143), .C(Rst_n), .D(n41), .Z(n3) );
  ND2M1P U77 ( .A(n64), .B(n10), .Z(n69) );
  OAI211M1P U78 ( .A(n146), .B(n145), .C(Rst_n), .D(n144), .Z(n375) );
  OAI211M1P U79 ( .A(n109), .B(n145), .C(Rst_n), .D(n144), .Z(n141) );
  AOI22M1P U80 ( .A(\Queue[3][0] ), .B(n51), .C(n374), .D(\Queue[4][0] ), .Z(
        n6) );
  OAI21M1P U81 ( .A(n149), .B(n377), .C(n6), .Z(n514) );
  OA21M1P U82 ( .A(n146), .B(n143), .C(n41), .Z(n7) );
  OAI21M1P U83 ( .A(n149), .B(n50), .C(n9), .Z(n482) );
  OAI21M1P U84 ( .A(n167), .B(n50), .C(n118), .Z(n491) );
  OAI21M1P U85 ( .A(n165), .B(n50), .C(n117), .Z(n490) );
  OAI21M1P U86 ( .A(n163), .B(n50), .C(n116), .Z(n489) );
  OAI21M1P U87 ( .A(n161), .B(n50), .C(n115), .Z(n488) );
  OAI21M1P U88 ( .A(n159), .B(n50), .C(n114), .Z(n487) );
  OAI21M1P U89 ( .A(n157), .B(n50), .C(n113), .Z(n486) );
  OAI21M1P U90 ( .A(n155), .B(n50), .C(n112), .Z(n485) );
  OAI21M1P U91 ( .A(n153), .B(n50), .C(n111), .Z(n484) );
  OAI21M1P U92 ( .A(n151), .B(n50), .C(n110), .Z(n483) );
  OA21M1P U93 ( .A(n145), .B(n109), .C(Rst_n), .Z(n8) );
  AOI22M1P U94 ( .A(\Queue[2][0] ), .B(n48), .C(\Queue[3][0] ), .D(n140), .Z(
        n9) );
  OA21M1P U95 ( .A(n109), .B(n143), .C(n41), .Z(n10) );
  AOI22M1P U96 ( .A(n68), .B(\Queue[2][16] ), .C(\Queue[1][16] ), .D(n43), .Z(
        n11) );
  OAI21M1P U97 ( .A(n44), .B(n181), .C(n11), .Z(n434) );
  AOI22M1P U98 ( .A(n68), .B(\Queue[2][31] ), .C(\Queue[1][31] ), .D(n42), .Z(
        n12) );
  OAI21M1P U99 ( .A(n45), .B(n378), .C(n12), .Z(n449) );
  AOI22M1P U100 ( .A(n68), .B(\Queue[2][8] ), .C(\Queue[1][8] ), .D(n42), .Z(
        n13) );
  OAI21M1P U101 ( .A(n44), .B(n165), .C(n13), .Z(n426) );
  AOI22M1P U102 ( .A(n68), .B(\Queue[2][30] ), .C(\Queue[1][30] ), .D(n42), 
        .Z(n14) );
  OAI21M1P U103 ( .A(n45), .B(n373), .C(n14), .Z(n448) );
  AOI22M1P U104 ( .A(n68), .B(\Queue[2][29] ), .C(\Queue[1][29] ), .D(n42), 
        .Z(n15) );
  OAI21M1P U105 ( .A(n45), .B(n207), .C(n15), .Z(n447) );
  AOI22M1P U106 ( .A(n68), .B(\Queue[2][15] ), .C(\Queue[1][15] ), .D(n43), 
        .Z(n16) );
  OAI21M1P U107 ( .A(n44), .B(n179), .C(n16), .Z(n433) );
  AOI22M1P U108 ( .A(n68), .B(\Queue[2][4] ), .C(\Queue[1][4] ), .D(n42), .Z(
        n17) );
  OAI21M1P U109 ( .A(n45), .B(n157), .C(n17), .Z(n422) );
  AOI22M1P U110 ( .A(n68), .B(\Queue[2][28] ), .C(\Queue[1][28] ), .D(n42), 
        .Z(n18) );
  OAI21M1P U111 ( .A(n45), .B(n205), .C(n18), .Z(n446) );
  AOI22M1P U112 ( .A(n68), .B(\Queue[2][27] ), .C(\Queue[1][27] ), .D(n42), 
        .Z(n19) );
  OAI21M1P U113 ( .A(n45), .B(n203), .C(n19), .Z(n445) );
  AOI22M1P U114 ( .A(n68), .B(\Queue[2][14] ), .C(\Queue[1][14] ), .D(n43), 
        .Z(n20) );
  OAI21M1P U115 ( .A(n44), .B(n177), .C(n20), .Z(n432) );
  AOI22M1P U116 ( .A(n68), .B(\Queue[2][23] ), .C(\Queue[1][23] ), .D(n43), 
        .Z(n21) );
  OAI21M1P U117 ( .A(n45), .B(n195), .C(n21), .Z(n441) );
  AOI22M1P U118 ( .A(n68), .B(\Queue[2][26] ), .C(\Queue[1][26] ), .D(n43), 
        .Z(n22) );
  OAI21M1P U119 ( .A(n45), .B(n201), .C(n22), .Z(n444) );
  AOI22M1P U120 ( .A(n68), .B(\Queue[2][2] ), .C(\Queue[1][2] ), .D(n42), .Z(
        n23) );
  OAI21M1P U121 ( .A(n44), .B(n153), .C(n23), .Z(n420) );
  AOI22M1P U122 ( .A(n68), .B(\Queue[2][13] ), .C(\Queue[1][13] ), .D(n43), 
        .Z(n24) );
  OAI21M1P U123 ( .A(n44), .B(n175), .C(n24), .Z(n431) );
  AOI22M1P U124 ( .A(n68), .B(\Queue[2][12] ), .C(\Queue[1][12] ), .D(n43), 
        .Z(n25) );
  OAI21M1P U125 ( .A(n44), .B(n173), .C(n25), .Z(n430) );
  AOI22M1P U126 ( .A(n68), .B(\Queue[2][24] ), .C(\Queue[1][24] ), .D(n43), 
        .Z(n26) );
  OAI21M1P U127 ( .A(n44), .B(n197), .C(n26), .Z(n442) );
  AOI22M1P U128 ( .A(n68), .B(\Queue[2][22] ), .C(\Queue[1][22] ), .D(n43), 
        .Z(n27) );
  OAI21M1P U129 ( .A(n45), .B(n193), .C(n27), .Z(n440) );
  AOI22M1P U130 ( .A(n68), .B(\Queue[2][6] ), .C(\Queue[1][6] ), .D(n42), .Z(
        n28) );
  OAI21M1P U131 ( .A(n45), .B(n161), .C(n28), .Z(n424) );
  AOI22M1P U132 ( .A(n68), .B(\Queue[2][21] ), .C(\Queue[1][21] ), .D(n43), 
        .Z(n29) );
  OAI21M1P U133 ( .A(n44), .B(n191), .C(n29), .Z(n439) );
  AOI22M1P U134 ( .A(n68), .B(\Queue[2][11] ), .C(\Queue[1][11] ), .D(n43), 
        .Z(n30) );
  OAI21M1P U135 ( .A(n44), .B(n171), .C(n30), .Z(n429) );
  AOI22M1P U136 ( .A(n68), .B(\Queue[2][10] ), .C(\Queue[1][10] ), .D(n43), 
        .Z(n31) );
  OAI21M1P U137 ( .A(n45), .B(n169), .C(n31), .Z(n428) );
  AOI22M1P U138 ( .A(n68), .B(\Queue[2][20] ), .C(\Queue[1][20] ), .D(n43), 
        .Z(n32) );
  OAI21M1P U139 ( .A(n44), .B(n189), .C(n32), .Z(n438) );
  AOI22M1P U140 ( .A(n68), .B(\Queue[2][19] ), .C(\Queue[1][19] ), .D(n43), 
        .Z(n33) );
  OAI21M1P U141 ( .A(n44), .B(n187), .C(n33), .Z(n437) );
  AOI22M1P U142 ( .A(n68), .B(\Queue[2][25] ), .C(\Queue[1][25] ), .D(n43), 
        .Z(n34) );
  OAI21M1P U143 ( .A(n45), .B(n199), .C(n34), .Z(n443) );
  AOI22M1P U144 ( .A(n68), .B(\Queue[2][3] ), .C(\Queue[1][3] ), .D(n42), .Z(
        n35) );
  OAI21M1P U145 ( .A(n69), .B(n155), .C(n35), .Z(n421) );
  AOI22M1P U146 ( .A(n68), .B(\Queue[2][18] ), .C(\Queue[1][18] ), .D(n43), 
        .Z(n36) );
  OAI21M1P U147 ( .A(n44), .B(n185), .C(n36), .Z(n436) );
  AOI22M1P U148 ( .A(n68), .B(\Queue[2][9] ), .C(\Queue[1][9] ), .D(n43), .Z(
        n37) );
  OAI21M1P U149 ( .A(n69), .B(n167), .C(n37), .Z(n427) );
  AOI22M1P U150 ( .A(n68), .B(\Queue[2][17] ), .C(\Queue[1][17] ), .D(n43), 
        .Z(n38) );
  OAI21M1P U151 ( .A(n44), .B(n183), .C(n38), .Z(n435) );
  AOI22M1P U152 ( .A(n68), .B(\Queue[2][5] ), .C(\Queue[1][5] ), .D(n42), .Z(
        n39) );
  OAI21M1P U153 ( .A(n69), .B(n159), .C(n39), .Z(n423) );
  AOI22M1P U154 ( .A(n68), .B(\Queue[2][7] ), .C(\Queue[1][7] ), .D(n42), .Z(
        n40) );
  OAI21M1P U155 ( .A(n69), .B(n163), .C(n40), .Z(n425) );
  NR2M1P U156 ( .A(n143), .B(n41), .Z(n380) );
  NR2M1P U157 ( .A(n58), .B(n380), .Z(n379) );
  AOI22CDNM1P U158 ( .A(n379), .B(n63), .C(n379), .D(n63), .Z(n382) );
  N1M1P U159 ( .A(n380), .Z(n57) );
  AOI22M1P U160 ( .A(Count[0]), .B(n145), .C(n57), .D(n63), .Z(n54) );
  AOI22CDNM1P U161 ( .A(Count[1]), .B(n54), .C(n54), .D(Count[1]), .Z(n383) );
  ND3M1P U162 ( .A(n63), .B(n59), .C(n62), .Z(n70) );
  ND2M1P U163 ( .A(Count[1]), .B(Read_Ack), .Z(n53) );
  OAI211M1P U164 ( .A(Count[1]), .B(n145), .C(n54), .D(n53), .Z(n55) );
  AOI22M1P U165 ( .A(n58), .B(n146), .C(Count[2]), .D(n55), .Z(n56) );
  OAI21M1P U166 ( .A(n70), .B(n57), .C(n56), .Z(n384) );
  AOI22CDNM1P U167 ( .A(n60), .B(n378), .C(\Queue[4][31] ), .D(n60), .Z(n385)
         );
  AOI22CDNM1P U168 ( .A(n60), .B(n149), .C(\Queue[4][0] ), .D(n60), .Z(n386)
         );
  AOI22CDNM1P U169 ( .A(n60), .B(n151), .C(\Queue[4][1] ), .D(n60), .Z(n387)
         );
  AOI22CDNM1P U170 ( .A(n60), .B(n153), .C(\Queue[4][2] ), .D(n60), .Z(n388)
         );
  AOI22CDNM1P U171 ( .A(n60), .B(n155), .C(\Queue[4][3] ), .D(n60), .Z(n389)
         );
  AOI22CDNM1P U172 ( .A(n60), .B(n157), .C(\Queue[4][4] ), .D(n60), .Z(n390)
         );
  AOI22CDNM1P U173 ( .A(n60), .B(n159), .C(\Queue[4][5] ), .D(n60), .Z(n391)
         );
  AOI22CDNM1P U174 ( .A(n60), .B(n161), .C(\Queue[4][6] ), .D(n60), .Z(n392)
         );
  AOI22CDNM1P U175 ( .A(n60), .B(n163), .C(\Queue[4][7] ), .D(n60), .Z(n393)
         );
  AOI22CDNM1P U176 ( .A(n60), .B(n165), .C(\Queue[4][8] ), .D(n60), .Z(n394)
         );
  AOI22CDNM1P U177 ( .A(n60), .B(n167), .C(\Queue[4][9] ), .D(n60), .Z(n395)
         );
  AOI22CDNM1P U178 ( .A(n60), .B(n169), .C(\Queue[4][10] ), .D(n60), .Z(n396)
         );
  AOI22CDNM1P U179 ( .A(n60), .B(n171), .C(\Queue[4][11] ), .D(n60), .Z(n397)
         );
  AOI22CDNM1P U180 ( .A(n60), .B(n173), .C(\Queue[4][12] ), .D(n60), .Z(n398)
         );
  AOI22CDNM1P U181 ( .A(n60), .B(n175), .C(\Queue[4][13] ), .D(n60), .Z(n399)
         );
  AOI22CDNM1P U182 ( .A(n60), .B(n177), .C(\Queue[4][14] ), .D(n60), .Z(n400)
         );
  AOI22CDNM1P U183 ( .A(n60), .B(n179), .C(\Queue[4][15] ), .D(n60), .Z(n401)
         );
  AOI22CDNM1P U184 ( .A(n60), .B(n181), .C(\Queue[4][16] ), .D(n60), .Z(n402)
         );
  AOI22CDNM1P U185 ( .A(n60), .B(n183), .C(\Queue[4][17] ), .D(n60), .Z(n403)
         );
  AOI22CDNM1P U186 ( .A(n60), .B(n185), .C(\Queue[4][18] ), .D(n60), .Z(n404)
         );
  AOI22CDNM1P U187 ( .A(n60), .B(n187), .C(\Queue[4][19] ), .D(n60), .Z(n405)
         );
  AOI22CDNM1P U188 ( .A(n60), .B(n189), .C(\Queue[4][20] ), .D(n60), .Z(n406)
         );
  AOI22CDNM1P U189 ( .A(n60), .B(n191), .C(\Queue[4][21] ), .D(n60), .Z(n407)
         );
  AOI22CDNM1P U190 ( .A(n60), .B(n193), .C(\Queue[4][22] ), .D(n60), .Z(n408)
         );
  AOI22CDNM1P U191 ( .A(n60), .B(n195), .C(\Queue[4][23] ), .D(n60), .Z(n409)
         );
  AOI22CDNM1P U192 ( .A(n60), .B(n197), .C(\Queue[4][24] ), .D(n60), .Z(n410)
         );
  AOI22CDNM1P U193 ( .A(n60), .B(n199), .C(\Queue[4][25] ), .D(n60), .Z(n411)
         );
  AOI22CDNM1P U194 ( .A(n60), .B(n201), .C(\Queue[4][26] ), .D(n60), .Z(n412)
         );
  AOI22CDNM1P U195 ( .A(n60), .B(n203), .C(\Queue[4][27] ), .D(n60), .Z(n413)
         );
  AOI22CDNM1P U196 ( .A(n60), .B(n205), .C(\Queue[4][28] ), .D(n60), .Z(n414)
         );
  AOI22CDNM1P U197 ( .A(n60), .B(n207), .C(\Queue[4][29] ), .D(n60), .Z(n415)
         );
  AOI22CDNM1P U198 ( .A(n60), .B(n373), .C(\Queue[4][30] ), .D(n60), .Z(n416)
         );
  OAI22CDNM1P U199 ( .A(n145), .B(n61), .C(n379), .D(Full), .Z(n417) );
  OAI21M1P U200 ( .A(n41), .B(Read_Ack), .C(n64), .Z(n67) );
  AOI22M1P U201 ( .A(n68), .B(\Queue[2][1] ), .C(\Queue[1][1] ), .D(n42), .Z(
        n66) );
  OAI21M1P U202 ( .A(n45), .B(n151), .C(n66), .Z(n419) );
  AOI22M1P U203 ( .A(\Queue[1][0] ), .B(n105), .C(n104), .D(Packet_Out[0]), 
        .Z(n73) );
  OAI21M1P U204 ( .A(n149), .B(n46), .C(n73), .Z(n450) );
  AOI22M1P U205 ( .A(\Queue[1][1] ), .B(n105), .C(n104), .D(Packet_Out[1]), 
        .Z(n74) );
  OAI21M1P U206 ( .A(n151), .B(n46), .C(n74), .Z(n451) );
  AOI22M1P U207 ( .A(\Queue[1][2] ), .B(n105), .C(n104), .D(Packet_Out[2]), 
        .Z(n75) );
  OAI21M1P U208 ( .A(n153), .B(n46), .C(n75), .Z(n452) );
  AOI22M1P U209 ( .A(\Queue[1][3] ), .B(n105), .C(n104), .D(Packet_Out[3]), 
        .Z(n76) );
  OAI21M1P U210 ( .A(n155), .B(n46), .C(n76), .Z(n453) );
  AOI22M1P U211 ( .A(\Queue[1][4] ), .B(n105), .C(n104), .D(Packet_Out[4]), 
        .Z(n77) );
  OAI21M1P U212 ( .A(n157), .B(n46), .C(n77), .Z(n454) );
  AOI22M1P U213 ( .A(\Queue[1][5] ), .B(n105), .C(n104), .D(Packet_Out[5]), 
        .Z(n78) );
  OAI21M1P U214 ( .A(n159), .B(n46), .C(n78), .Z(n455) );
  AOI22M1P U215 ( .A(\Queue[1][6] ), .B(n105), .C(n104), .D(Packet_Out[6]), 
        .Z(n79) );
  OAI21M1P U216 ( .A(n161), .B(n46), .C(n79), .Z(n456) );
  AOI22M1P U217 ( .A(\Queue[1][7] ), .B(n105), .C(n104), .D(Packet_Out[7]), 
        .Z(n80) );
  OAI21M1P U218 ( .A(n163), .B(n46), .C(n80), .Z(n457) );
  AOI22M1P U219 ( .A(\Queue[1][8] ), .B(n105), .C(n104), .D(Packet_Out[8]), 
        .Z(n81) );
  OAI21M1P U220 ( .A(n165), .B(n46), .C(n81), .Z(n458) );
  AOI22M1P U221 ( .A(\Queue[1][9] ), .B(n105), .C(n104), .D(Packet_Out[9]), 
        .Z(n82) );
  OAI21M1P U222 ( .A(n167), .B(n46), .C(n82), .Z(n459) );
  AOI22M1P U223 ( .A(\Queue[1][10] ), .B(n105), .C(n104), .D(Packet_Out[10]), 
        .Z(n83) );
  OAI21M1P U224 ( .A(n169), .B(n47), .C(n83), .Z(n460) );
  AOI22M1P U225 ( .A(\Queue[1][11] ), .B(n105), .C(n104), .D(Packet_Out[11]), 
        .Z(n84) );
  OAI21M1P U226 ( .A(n171), .B(n47), .C(n84), .Z(n461) );
  AOI22M1P U227 ( .A(\Queue[1][12] ), .B(n105), .C(n104), .D(Packet_Out[12]), 
        .Z(n85) );
  OAI21M1P U228 ( .A(n173), .B(n47), .C(n85), .Z(n462) );
  AOI22M1P U229 ( .A(\Queue[1][13] ), .B(n105), .C(n104), .D(Packet_Out[13]), 
        .Z(n86) );
  OAI21M1P U230 ( .A(n175), .B(n47), .C(n86), .Z(n463) );
  AOI22M1P U231 ( .A(\Queue[1][14] ), .B(n105), .C(n104), .D(Packet_Out[14]), 
        .Z(n87) );
  OAI21M1P U232 ( .A(n177), .B(n47), .C(n87), .Z(n464) );
  AOI22M1P U233 ( .A(\Queue[1][15] ), .B(n105), .C(n104), .D(Packet_Out[15]), 
        .Z(n88) );
  OAI21M1P U234 ( .A(n179), .B(n47), .C(n88), .Z(n465) );
  AOI22M1P U235 ( .A(\Queue[1][16] ), .B(n105), .C(n104), .D(Packet_Out[16]), 
        .Z(n89) );
  OAI21M1P U236 ( .A(n181), .B(n47), .C(n89), .Z(n466) );
  AOI22M1P U237 ( .A(\Queue[1][17] ), .B(n105), .C(n104), .D(Packet_Out[17]), 
        .Z(n90) );
  OAI21M1P U238 ( .A(n183), .B(n47), .C(n90), .Z(n467) );
  AOI22M1P U239 ( .A(\Queue[1][18] ), .B(n105), .C(n104), .D(Packet_Out[18]), 
        .Z(n91) );
  OAI21M1P U240 ( .A(n185), .B(n47), .C(n91), .Z(n468) );
  AOI22M1P U241 ( .A(\Queue[1][19] ), .B(n105), .C(n104), .D(Packet_Out[19]), 
        .Z(n92) );
  OAI21M1P U242 ( .A(n187), .B(n47), .C(n92), .Z(n469) );
  AOI22M1P U243 ( .A(\Queue[1][20] ), .B(n105), .C(n104), .D(Packet_Out[20]), 
        .Z(n93) );
  OAI21M1P U244 ( .A(n189), .B(n47), .C(n93), .Z(n470) );
  AOI22M1P U245 ( .A(\Queue[1][21] ), .B(n105), .C(n104), .D(Packet_Out[21]), 
        .Z(n94) );
  OAI21M1P U246 ( .A(n191), .B(n47), .C(n94), .Z(n471) );
  AOI22M1P U247 ( .A(\Queue[1][22] ), .B(n105), .C(n104), .D(Packet_Out[22]), 
        .Z(n95) );
  OAI21M1P U248 ( .A(n193), .B(n47), .C(n95), .Z(n472) );
  AOI22M1P U249 ( .A(\Queue[1][23] ), .B(n105), .C(n104), .D(Packet_Out[23]), 
        .Z(n96) );
  OAI21M1P U250 ( .A(n195), .B(n47), .C(n96), .Z(n473) );
  AOI22M1P U251 ( .A(\Queue[1][24] ), .B(n105), .C(n104), .D(Packet_Out[24]), 
        .Z(n97) );
  OAI21M1P U252 ( .A(n197), .B(n47), .C(n97), .Z(n474) );
  AOI22M1P U253 ( .A(\Queue[1][25] ), .B(n105), .C(n104), .D(Packet_Out[25]), 
        .Z(n98) );
  OAI21M1P U254 ( .A(n199), .B(n47), .C(n98), .Z(n475) );
  AOI22M1P U255 ( .A(\Queue[1][26] ), .B(n105), .C(n104), .D(Packet_Out[26]), 
        .Z(n99) );
  OAI21M1P U256 ( .A(n201), .B(n47), .C(n99), .Z(n476) );
  AOI22M1P U257 ( .A(\Queue[1][27] ), .B(n105), .C(n104), .D(Packet_Out[27]), 
        .Z(n100) );
  OAI21M1P U258 ( .A(n203), .B(n47), .C(n100), .Z(n477) );
  AOI22M1P U259 ( .A(\Queue[1][28] ), .B(n105), .C(n104), .D(Packet_Out[28]), 
        .Z(n101) );
  OAI21M1P U260 ( .A(n205), .B(n47), .C(n101), .Z(n478) );
  AOI22M1P U261 ( .A(\Queue[1][29] ), .B(n105), .C(n104), .D(Packet_Out[29]), 
        .Z(n102) );
  OAI21M1P U262 ( .A(n207), .B(n47), .C(n102), .Z(n479) );
  AOI22M1P U263 ( .A(\Queue[1][30] ), .B(n105), .C(n104), .D(Packet_Out[30]), 
        .Z(n103) );
  OAI21M1P U264 ( .A(n373), .B(n46), .C(n103), .Z(n480) );
  AOI22M1P U265 ( .A(\Queue[1][31] ), .B(n105), .C(n104), .D(Packet_Out[31]), 
        .Z(n106) );
  OAI21M1P U266 ( .A(n378), .B(n47), .C(n106), .Z(n481) );
  ND2M1P U267 ( .A(n108), .B(n143), .Z(n144) );
  AOI22M1P U268 ( .A(\Queue[2][2] ), .B(n48), .C(n140), .D(\Queue[3][2] ), .Z(
        n111) );
  AOI22M1P U269 ( .A(\Queue[2][3] ), .B(n48), .C(n140), .D(\Queue[3][3] ), .Z(
        n112) );
  AOI22M1P U270 ( .A(\Queue[2][4] ), .B(n48), .C(n140), .D(\Queue[3][4] ), .Z(
        n113) );
  AOI22M1P U271 ( .A(\Queue[2][5] ), .B(n48), .C(n140), .D(\Queue[3][5] ), .Z(
        n114) );
  AOI22M1P U272 ( .A(\Queue[2][6] ), .B(n48), .C(n140), .D(\Queue[3][6] ), .Z(
        n115) );
  AOI22M1P U273 ( .A(\Queue[2][7] ), .B(n48), .C(n140), .D(\Queue[3][7] ), .Z(
        n116) );
  AOI22M1P U274 ( .A(\Queue[2][8] ), .B(n48), .C(n140), .D(\Queue[3][8] ), .Z(
        n117) );
  AOI22M1P U275 ( .A(\Queue[2][9] ), .B(n48), .C(n140), .D(\Queue[3][9] ), .Z(
        n118) );
  AOI22M1P U276 ( .A(\Queue[2][10] ), .B(n48), .C(n140), .D(\Queue[3][10] ), 
        .Z(n119) );
  OAI21M1P U277 ( .A(n169), .B(n50), .C(n119), .Z(n492) );
  AOI22M1P U278 ( .A(\Queue[2][11] ), .B(n48), .C(n140), .D(\Queue[3][11] ), 
        .Z(n120) );
  OAI21M1P U279 ( .A(n171), .B(n50), .C(n120), .Z(n493) );
  AOI22M1P U280 ( .A(\Queue[2][12] ), .B(n48), .C(n140), .D(\Queue[3][12] ), 
        .Z(n121) );
  OAI21M1P U281 ( .A(n173), .B(n50), .C(n121), .Z(n494) );
  AOI22M1P U282 ( .A(\Queue[2][13] ), .B(n48), .C(n140), .D(\Queue[3][13] ), 
        .Z(n122) );
  OAI21M1P U283 ( .A(n175), .B(n50), .C(n122), .Z(n495) );
  AOI22M1P U284 ( .A(\Queue[2][14] ), .B(n48), .C(n140), .D(\Queue[3][14] ), 
        .Z(n123) );
  OAI21M1P U285 ( .A(n177), .B(n50), .C(n123), .Z(n496) );
  AOI22M1P U286 ( .A(\Queue[2][15] ), .B(n48), .C(n140), .D(\Queue[3][15] ), 
        .Z(n124) );
  OAI21M1P U287 ( .A(n179), .B(n50), .C(n124), .Z(n497) );
  AOI22M1P U288 ( .A(\Queue[2][16] ), .B(n48), .C(n140), .D(\Queue[3][16] ), 
        .Z(n125) );
  OAI21M1P U289 ( .A(n181), .B(n50), .C(n125), .Z(n498) );
  AOI22M1P U290 ( .A(\Queue[2][17] ), .B(n48), .C(n140), .D(\Queue[3][17] ), 
        .Z(n126) );
  OAI21M1P U291 ( .A(n183), .B(n50), .C(n126), .Z(n499) );
  AOI22M1P U292 ( .A(\Queue[2][18] ), .B(n48), .C(n140), .D(\Queue[3][18] ), 
        .Z(n127) );
  OAI21M1P U293 ( .A(n185), .B(n50), .C(n127), .Z(n500) );
  AOI22M1P U294 ( .A(\Queue[2][19] ), .B(n48), .C(n140), .D(\Queue[3][19] ), 
        .Z(n128) );
  OAI21M1P U295 ( .A(n187), .B(n50), .C(n128), .Z(n501) );
  AOI22M1P U296 ( .A(\Queue[2][20] ), .B(n49), .C(n140), .D(\Queue[3][20] ), 
        .Z(n129) );
  OAI21M1P U297 ( .A(n189), .B(n50), .C(n129), .Z(n502) );
  AOI22M1P U298 ( .A(\Queue[2][21] ), .B(n49), .C(n140), .D(\Queue[3][21] ), 
        .Z(n130) );
  OAI21M1P U299 ( .A(n191), .B(n50), .C(n130), .Z(n503) );
  AOI22M1P U300 ( .A(\Queue[2][22] ), .B(n49), .C(n140), .D(\Queue[3][22] ), 
        .Z(n131) );
  OAI21M1P U301 ( .A(n193), .B(n50), .C(n131), .Z(n504) );
  AOI22M1P U302 ( .A(\Queue[2][23] ), .B(n49), .C(n140), .D(\Queue[3][23] ), 
        .Z(n132) );
  OAI21M1P U303 ( .A(n195), .B(n50), .C(n132), .Z(n505) );
  AOI22M1P U304 ( .A(\Queue[2][24] ), .B(n49), .C(n140), .D(\Queue[3][24] ), 
        .Z(n133) );
  OAI21M1P U305 ( .A(n197), .B(n50), .C(n133), .Z(n506) );
  AOI22M1P U306 ( .A(\Queue[2][25] ), .B(n49), .C(n140), .D(\Queue[3][25] ), 
        .Z(n134) );
  OAI21M1P U307 ( .A(n199), .B(n50), .C(n134), .Z(n507) );
  AOI22M1P U308 ( .A(\Queue[2][26] ), .B(n49), .C(n140), .D(\Queue[3][26] ), 
        .Z(n135) );
  OAI21M1P U309 ( .A(n201), .B(n50), .C(n135), .Z(n508) );
  AOI22M1P U310 ( .A(\Queue[2][27] ), .B(n49), .C(n140), .D(\Queue[3][27] ), 
        .Z(n136) );
  OAI21M1P U311 ( .A(n203), .B(n50), .C(n136), .Z(n509) );
  AOI22M1P U312 ( .A(\Queue[2][28] ), .B(n49), .C(n140), .D(\Queue[3][28] ), 
        .Z(n137) );
  OAI21M1P U313 ( .A(n205), .B(n50), .C(n137), .Z(n510) );
  AOI22M1P U314 ( .A(\Queue[2][29] ), .B(n49), .C(n140), .D(\Queue[3][29] ), 
        .Z(n138) );
  OAI21M1P U315 ( .A(n207), .B(n50), .C(n138), .Z(n511) );
  AOI22M1P U316 ( .A(\Queue[2][30] ), .B(n48), .C(n140), .D(\Queue[3][30] ), 
        .Z(n139) );
  OAI21M1P U317 ( .A(n373), .B(n50), .C(n139), .Z(n512) );
  AOI22M1P U318 ( .A(\Queue[2][31] ), .B(n49), .C(n140), .D(\Queue[3][31] ), 
        .Z(n142) );
  OAI21M1P U319 ( .A(n378), .B(n50), .C(n142), .Z(n513) );
  AOI22M1P U320 ( .A(\Queue[3][1] ), .B(n51), .C(n374), .D(\Queue[4][1] ), .Z(
        n150) );
  OAI21M1P U321 ( .A(n151), .B(n377), .C(n150), .Z(n515) );
  AOI22M1P U322 ( .A(\Queue[3][2] ), .B(n51), .C(n374), .D(\Queue[4][2] ), .Z(
        n152) );
  OAI21M1P U323 ( .A(n153), .B(n377), .C(n152), .Z(n516) );
  AOI22M1P U324 ( .A(\Queue[3][3] ), .B(n51), .C(n374), .D(\Queue[4][3] ), .Z(
        n154) );
  OAI21M1P U325 ( .A(n155), .B(n377), .C(n154), .Z(n517) );
  AOI22M1P U326 ( .A(\Queue[3][4] ), .B(n51), .C(n374), .D(\Queue[4][4] ), .Z(
        n156) );
  OAI21M1P U327 ( .A(n157), .B(n377), .C(n156), .Z(n518) );
  AOI22M1P U328 ( .A(\Queue[3][5] ), .B(n51), .C(n374), .D(\Queue[4][5] ), .Z(
        n158) );
  OAI21M1P U329 ( .A(n159), .B(n377), .C(n158), .Z(n519) );
  AOI22M1P U330 ( .A(\Queue[3][6] ), .B(n51), .C(n374), .D(\Queue[4][6] ), .Z(
        n160) );
  OAI21M1P U331 ( .A(n161), .B(n377), .C(n160), .Z(n520) );
  AOI22M1P U332 ( .A(\Queue[3][7] ), .B(n51), .C(n374), .D(\Queue[4][7] ), .Z(
        n162) );
  OAI21M1P U333 ( .A(n163), .B(n377), .C(n162), .Z(n521) );
  AOI22M1P U334 ( .A(\Queue[3][8] ), .B(n51), .C(n374), .D(\Queue[4][8] ), .Z(
        n164) );
  OAI21M1P U335 ( .A(n165), .B(n377), .C(n164), .Z(n522) );
  AOI22M1P U336 ( .A(\Queue[3][9] ), .B(n51), .C(n374), .D(\Queue[4][9] ), .Z(
        n166) );
  OAI21M1P U337 ( .A(n167), .B(n377), .C(n166), .Z(n523) );
  AOI22M1P U338 ( .A(\Queue[3][10] ), .B(n51), .C(n374), .D(\Queue[4][10] ), 
        .Z(n168) );
  OAI21M1P U339 ( .A(n169), .B(n377), .C(n168), .Z(n524) );
  AOI22M1P U340 ( .A(\Queue[3][11] ), .B(n51), .C(n374), .D(\Queue[4][11] ), 
        .Z(n170) );
  OAI21M1P U341 ( .A(n171), .B(n377), .C(n170), .Z(n525) );
  AOI22M1P U342 ( .A(\Queue[3][12] ), .B(n51), .C(n374), .D(\Queue[4][12] ), 
        .Z(n172) );
  OAI21M1P U343 ( .A(n173), .B(n377), .C(n172), .Z(n526) );
  AOI22M1P U344 ( .A(\Queue[3][13] ), .B(n51), .C(n374), .D(\Queue[4][13] ), 
        .Z(n174) );
  OAI21M1P U345 ( .A(n175), .B(n377), .C(n174), .Z(n527) );
  AOI22M1P U346 ( .A(\Queue[3][14] ), .B(n51), .C(n374), .D(\Queue[4][14] ), 
        .Z(n176) );
  OAI21M1P U347 ( .A(n177), .B(n377), .C(n176), .Z(n528) );
  AOI22M1P U348 ( .A(\Queue[3][15] ), .B(n51), .C(n374), .D(\Queue[4][15] ), 
        .Z(n178) );
  OAI21M1P U349 ( .A(n179), .B(n377), .C(n178), .Z(n529) );
  AOI22M1P U350 ( .A(\Queue[3][16] ), .B(n51), .C(n374), .D(\Queue[4][16] ), 
        .Z(n180) );
  OAI21M1P U351 ( .A(n181), .B(n377), .C(n180), .Z(n530) );
  AOI22M1P U352 ( .A(\Queue[3][17] ), .B(n51), .C(n374), .D(\Queue[4][17] ), 
        .Z(n182) );
  OAI21M1P U353 ( .A(n183), .B(n377), .C(n182), .Z(n531) );
  AOI22M1P U354 ( .A(\Queue[3][18] ), .B(n51), .C(n374), .D(\Queue[4][18] ), 
        .Z(n184) );
  OAI21M1P U355 ( .A(n185), .B(n377), .C(n184), .Z(n532) );
  AOI22M1P U356 ( .A(\Queue[3][19] ), .B(n51), .C(n374), .D(\Queue[4][19] ), 
        .Z(n186) );
  OAI21M1P U357 ( .A(n187), .B(n377), .C(n186), .Z(n533) );
  AOI22M1P U358 ( .A(\Queue[3][20] ), .B(n52), .C(n374), .D(\Queue[4][20] ), 
        .Z(n188) );
  OAI21M1P U359 ( .A(n189), .B(n377), .C(n188), .Z(n534) );
  AOI22M1P U360 ( .A(\Queue[3][21] ), .B(n52), .C(n374), .D(\Queue[4][21] ), 
        .Z(n190) );
  OAI21M1P U361 ( .A(n191), .B(n377), .C(n190), .Z(n535) );
  AOI22M1P U362 ( .A(\Queue[3][22] ), .B(n52), .C(n374), .D(\Queue[4][22] ), 
        .Z(n192) );
  OAI21M1P U363 ( .A(n193), .B(n377), .C(n192), .Z(n536) );
  AOI22M1P U364 ( .A(\Queue[3][23] ), .B(n52), .C(n374), .D(\Queue[4][23] ), 
        .Z(n194) );
  OAI21M1P U365 ( .A(n195), .B(n377), .C(n194), .Z(n537) );
  AOI22M1P U366 ( .A(\Queue[3][24] ), .B(n52), .C(n374), .D(\Queue[4][24] ), 
        .Z(n196) );
  OAI21M1P U367 ( .A(n197), .B(n377), .C(n196), .Z(n538) );
  AOI22M1P U368 ( .A(\Queue[3][25] ), .B(n52), .C(n374), .D(\Queue[4][25] ), 
        .Z(n198) );
  OAI21M1P U369 ( .A(n199), .B(n377), .C(n198), .Z(n539) );
  AOI22M1P U370 ( .A(\Queue[3][26] ), .B(n52), .C(n374), .D(\Queue[4][26] ), 
        .Z(n200) );
  OAI21M1P U371 ( .A(n201), .B(n377), .C(n200), .Z(n540) );
  AOI22M1P U372 ( .A(\Queue[3][27] ), .B(n52), .C(n374), .D(\Queue[4][27] ), 
        .Z(n202) );
  OAI21M1P U373 ( .A(n203), .B(n377), .C(n202), .Z(n541) );
  AOI22M1P U374 ( .A(\Queue[3][28] ), .B(n52), .C(n374), .D(\Queue[4][28] ), 
        .Z(n204) );
  OAI21M1P U375 ( .A(n205), .B(n377), .C(n204), .Z(n542) );
  AOI22M1P U376 ( .A(\Queue[3][29] ), .B(n52), .C(n374), .D(\Queue[4][29] ), 
        .Z(n206) );
  OAI21M1P U377 ( .A(n207), .B(n377), .C(n206), .Z(n543) );
  AOI22M1P U378 ( .A(\Queue[3][30] ), .B(n51), .C(n374), .D(\Queue[4][30] ), 
        .Z(n208) );
  OAI21M1P U379 ( .A(n373), .B(n377), .C(n208), .Z(n544) );
  AOI22M1P U380 ( .A(\Queue[3][31] ), .B(n52), .C(n374), .D(\Queue[4][31] ), 
        .Z(n376) );
  OAI21M1P U381 ( .A(n378), .B(n377), .C(n376), .Z(n545) );
  N1M1P U382 ( .A(n546), .Z(Empty) );
  AOI22M1P U383 ( .A(n381), .B(n380), .C(n379), .D(Empty), .Z(n547) );
endmodule


module Link_Control_2 ( Clk_r, Rst_n, Tx_Ready, Tx_Error, RxData_Valid, RxData, 
        Packet_From_Core, TxQueue_Write, RxQueue_Read, TxData_Valid, TxData, 
        Error_Ack, Core_Rcv_Ready, Packet_To_Core, RxQueue_Empty, TxQueue_Full
 );
  input [31:0] RxData;
  input [31:0] Packet_From_Core;
  output [31:0] TxData;
  output [31:0] Packet_To_Core;
  input Clk_r, Rst_n, Tx_Ready, Tx_Error, RxData_Valid, TxQueue_Write,
         RxQueue_Read;
  output TxData_Valid, Error_Ack, Core_Rcv_Ready, RxQueue_Empty, TxQueue_Full;
  wire   TxQueue_Read, TxQueue_Empty, RxQueue_Write, RxQueue_Full, N9, N16, n5,
         n6, n7, n8, n9;

  Packet_Queue_6 TxQueue ( .Clk_r(Clk_r), .Rst_n(Rst_n), .Packet_In(
        Packet_From_Core), .Read_Ack(TxQueue_Read), .Write_Ack(TxQueue_Write), 
        .Packet_Out(TxData), .Empty(TxQueue_Empty), .Full(TxQueue_Full) );
  Packet_Queue_5 RxQueue ( .Clk_r(Clk_r), .Rst_n(Rst_n), .Packet_In(RxData), 
        .Read_Ack(RxQueue_Read), .Write_Ack(RxQueue_Write), .Packet_Out(
        Packet_To_Core), .Empty(RxQueue_Empty), .Full(RxQueue_Full) );
  FD2QM1P Core_Rcv_Ready_reg ( .D(N9), .CP(Clk_r), .CD(Rst_n), .Q(
        Core_Rcv_Ready) );
  FD2QM1P TxQueue_Read_reg ( .D(N16), .CP(Clk_r), .CD(Rst_n), .Q(TxQueue_Read)
         );
  FD4QM1P RxQueue_Write_reg ( .D(n7), .CP(Clk_r), .SD(Rst_n), .Q(n6) );
  FD4QM1P TxData_Valid_reg ( .D(n9), .CP(Clk_r), .SD(Rst_n), .Q(n8) );
  N1M3P U3 ( .A(n6), .Z(RxQueue_Write) );
  NR2M1P U4 ( .A(n8), .B(Tx_Ready), .Z(N16) );
  NR2M1P U5 ( .A(RxData_Valid), .B(RxQueue_Full), .Z(n5) );
  OA21M1P U6 ( .A(Core_Rcv_Ready), .B(n5), .C(n6), .Z(N9) );
  N1M1P U7 ( .A(n8), .Z(TxData_Valid) );
  ND3M1P U8 ( .A(n6), .B(Core_Rcv_Ready), .C(RxData_Valid), .Z(n7) );
  AO21CNM1P U9 ( .A(n8), .B(TxQueue_Empty), .C(Tx_Ready), .Z(n9) );
endmodule


module Packet_Queue_7 ( Clk_r, Rst_n, Packet_In, Read_Ack, Write_Ack, 
        Packet_Out, Empty, Full );
  input [31:0] Packet_In;
  output [31:0] Packet_Out;
  input Clk_r, Rst_n, Read_Ack, Write_Ack;
  output Empty, Full;
  wire   \Queue[4][31] , \Queue[4][30] , \Queue[4][29] , \Queue[4][28] ,
         \Queue[4][27] , \Queue[4][26] , \Queue[4][25] , \Queue[4][24] ,
         \Queue[4][23] , \Queue[4][22] , \Queue[4][21] , \Queue[4][20] ,
         \Queue[4][19] , \Queue[4][18] , \Queue[4][17] , \Queue[4][16] ,
         \Queue[4][15] , \Queue[4][14] , \Queue[4][13] , \Queue[4][12] ,
         \Queue[4][11] , \Queue[4][10] , \Queue[4][9] , \Queue[4][8] ,
         \Queue[4][7] , \Queue[4][6] , \Queue[4][5] , \Queue[4][4] ,
         \Queue[4][3] , \Queue[4][2] , \Queue[4][1] , \Queue[4][0] ,
         \Queue[3][31] , \Queue[3][30] , \Queue[3][29] , \Queue[3][28] ,
         \Queue[3][27] , \Queue[3][26] , \Queue[3][25] , \Queue[3][24] ,
         \Queue[3][23] , \Queue[3][22] , \Queue[3][21] , \Queue[3][20] ,
         \Queue[3][19] , \Queue[3][18] , \Queue[3][17] , \Queue[3][16] ,
         \Queue[3][15] , \Queue[3][14] , \Queue[3][13] , \Queue[3][12] ,
         \Queue[3][11] , \Queue[3][10] , \Queue[3][9] , \Queue[3][8] ,
         \Queue[3][7] , \Queue[3][6] , \Queue[3][5] , \Queue[3][4] ,
         \Queue[3][3] , \Queue[3][2] , \Queue[3][1] , \Queue[3][0] ,
         \Queue[2][31] , \Queue[2][30] , \Queue[2][29] , \Queue[2][28] ,
         \Queue[2][27] , \Queue[2][26] , \Queue[2][25] , \Queue[2][24] ,
         \Queue[2][23] , \Queue[2][22] , \Queue[2][21] , \Queue[2][20] ,
         \Queue[2][19] , \Queue[2][18] , \Queue[2][17] , \Queue[2][16] ,
         \Queue[2][15] , \Queue[2][14] , \Queue[2][13] , \Queue[2][12] ,
         \Queue[2][11] , \Queue[2][10] , \Queue[2][9] , \Queue[2][8] ,
         \Queue[2][7] , \Queue[2][6] , \Queue[2][5] , \Queue[2][4] ,
         \Queue[2][3] , \Queue[2][2] , \Queue[2][1] , \Queue[2][0] ,
         \Queue[1][31] , \Queue[1][30] , \Queue[1][29] , \Queue[1][28] ,
         \Queue[1][27] , \Queue[1][26] , \Queue[1][25] , \Queue[1][24] ,
         \Queue[1][23] , \Queue[1][22] , \Queue[1][21] , \Queue[1][20] ,
         \Queue[1][19] , \Queue[1][18] , \Queue[1][17] , \Queue[1][16] ,
         \Queue[1][15] , \Queue[1][14] , \Queue[1][13] , \Queue[1][12] ,
         \Queue[1][11] , \Queue[1][10] , \Queue[1][9] , \Queue[1][8] ,
         \Queue[1][7] , \Queue[1][6] , \Queue[1][5] , \Queue[1][4] ,
         \Queue[1][3] , \Queue[1][2] , \Queue[1][1] , \Queue[1][0] , n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539;
  wire   [2:0] Count;

  FDN2QM1P \Count_reg[0]  ( .D(n374), .CPN(Clk_r), .CD(Rst_n), .Q(Count[0]) );
  FDN2QM1P \Count_reg[1]  ( .D(n375), .CPN(Clk_r), .CD(Rst_n), .Q(Count[1]) );
  FDN2QM1P \Count_reg[2]  ( .D(n376), .CPN(Clk_r), .CD(Rst_n), .Q(Count[2]) );
  FDN1QM1P \Queue_reg[4][30]  ( .D(n408), .CPN(Clk_r), .Q(\Queue[4][30] ) );
  FDN1QM1P \Queue_reg[3][30]  ( .D(n536), .CPN(Clk_r), .Q(\Queue[3][30] ) );
  FDN1QM1P \Queue_reg[2][30]  ( .D(n504), .CPN(Clk_r), .Q(\Queue[2][30] ) );
  FDN1QM1P \Queue_reg[4][29]  ( .D(n407), .CPN(Clk_r), .Q(\Queue[4][29] ) );
  FDN1QM1P \Queue_reg[3][29]  ( .D(n535), .CPN(Clk_r), .Q(\Queue[3][29] ) );
  FDN1QM1P \Queue_reg[2][29]  ( .D(n503), .CPN(Clk_r), .Q(\Queue[2][29] ) );
  FDN1QM1P \Queue_reg[4][28]  ( .D(n406), .CPN(Clk_r), .Q(\Queue[4][28] ) );
  FDN1QM1P \Queue_reg[3][28]  ( .D(n534), .CPN(Clk_r), .Q(\Queue[3][28] ) );
  FDN1QM1P \Queue_reg[2][28]  ( .D(n502), .CPN(Clk_r), .Q(\Queue[2][28] ) );
  FDN1QM1P \Queue_reg[4][27]  ( .D(n405), .CPN(Clk_r), .Q(\Queue[4][27] ) );
  FDN1QM1P \Queue_reg[3][27]  ( .D(n533), .CPN(Clk_r), .Q(\Queue[3][27] ) );
  FDN1QM1P \Queue_reg[2][27]  ( .D(n501), .CPN(Clk_r), .Q(\Queue[2][27] ) );
  FDN1QM1P \Queue_reg[4][26]  ( .D(n404), .CPN(Clk_r), .Q(\Queue[4][26] ) );
  FDN1QM1P \Queue_reg[3][26]  ( .D(n532), .CPN(Clk_r), .Q(\Queue[3][26] ) );
  FDN1QM1P \Queue_reg[2][26]  ( .D(n500), .CPN(Clk_r), .Q(\Queue[2][26] ) );
  FDN1QM1P \Queue_reg[4][25]  ( .D(n403), .CPN(Clk_r), .Q(\Queue[4][25] ) );
  FDN1QM1P \Queue_reg[3][25]  ( .D(n531), .CPN(Clk_r), .Q(\Queue[3][25] ) );
  FDN1QM1P \Queue_reg[2][25]  ( .D(n499), .CPN(Clk_r), .Q(\Queue[2][25] ) );
  FDN1QM1P \Queue_reg[4][24]  ( .D(n402), .CPN(Clk_r), .Q(\Queue[4][24] ) );
  FDN1QM1P \Queue_reg[3][24]  ( .D(n530), .CPN(Clk_r), .Q(\Queue[3][24] ) );
  FDN1QM1P \Queue_reg[2][24]  ( .D(n498), .CPN(Clk_r), .Q(\Queue[2][24] ) );
  FDN1QM1P \Queue_reg[4][23]  ( .D(n401), .CPN(Clk_r), .Q(\Queue[4][23] ) );
  FDN1QM1P \Queue_reg[3][23]  ( .D(n529), .CPN(Clk_r), .Q(\Queue[3][23] ) );
  FDN1QM1P \Queue_reg[2][23]  ( .D(n497), .CPN(Clk_r), .Q(\Queue[2][23] ) );
  FDN1QM1P \Queue_reg[4][22]  ( .D(n400), .CPN(Clk_r), .Q(\Queue[4][22] ) );
  FDN1QM1P \Queue_reg[3][22]  ( .D(n528), .CPN(Clk_r), .Q(\Queue[3][22] ) );
  FDN1QM1P \Queue_reg[2][22]  ( .D(n496), .CPN(Clk_r), .Q(\Queue[2][22] ) );
  FDN1QM1P \Queue_reg[4][21]  ( .D(n399), .CPN(Clk_r), .Q(\Queue[4][21] ) );
  FDN1QM1P \Queue_reg[3][21]  ( .D(n527), .CPN(Clk_r), .Q(\Queue[3][21] ) );
  FDN1QM1P \Queue_reg[2][21]  ( .D(n495), .CPN(Clk_r), .Q(\Queue[2][21] ) );
  FDN1QM1P \Queue_reg[4][20]  ( .D(n398), .CPN(Clk_r), .Q(\Queue[4][20] ) );
  FDN1QM1P \Queue_reg[3][20]  ( .D(n526), .CPN(Clk_r), .Q(\Queue[3][20] ) );
  FDN1QM1P \Queue_reg[2][20]  ( .D(n494), .CPN(Clk_r), .Q(\Queue[2][20] ) );
  FDN1QM1P \Queue_reg[4][19]  ( .D(n397), .CPN(Clk_r), .Q(\Queue[4][19] ) );
  FDN1QM1P \Queue_reg[3][19]  ( .D(n525), .CPN(Clk_r), .Q(\Queue[3][19] ) );
  FDN1QM1P \Queue_reg[2][19]  ( .D(n493), .CPN(Clk_r), .Q(\Queue[2][19] ) );
  FDN1QM1P \Queue_reg[4][18]  ( .D(n396), .CPN(Clk_r), .Q(\Queue[4][18] ) );
  FDN1QM1P \Queue_reg[3][18]  ( .D(n524), .CPN(Clk_r), .Q(\Queue[3][18] ) );
  FDN1QM1P \Queue_reg[2][18]  ( .D(n492), .CPN(Clk_r), .Q(\Queue[2][18] ) );
  FDN1QM1P \Queue_reg[4][17]  ( .D(n395), .CPN(Clk_r), .Q(\Queue[4][17] ) );
  FDN1QM1P \Queue_reg[3][17]  ( .D(n523), .CPN(Clk_r), .Q(\Queue[3][17] ) );
  FDN1QM1P \Queue_reg[2][17]  ( .D(n491), .CPN(Clk_r), .Q(\Queue[2][17] ) );
  FDN1QM1P \Queue_reg[4][16]  ( .D(n394), .CPN(Clk_r), .Q(\Queue[4][16] ) );
  FDN1QM1P \Queue_reg[3][16]  ( .D(n522), .CPN(Clk_r), .Q(\Queue[3][16] ) );
  FDN1QM1P \Queue_reg[2][16]  ( .D(n490), .CPN(Clk_r), .Q(\Queue[2][16] ) );
  FDN1QM1P \Queue_reg[4][15]  ( .D(n393), .CPN(Clk_r), .Q(\Queue[4][15] ) );
  FDN1QM1P \Queue_reg[3][15]  ( .D(n521), .CPN(Clk_r), .Q(\Queue[3][15] ) );
  FDN1QM1P \Queue_reg[2][15]  ( .D(n489), .CPN(Clk_r), .Q(\Queue[2][15] ) );
  FDN1QM1P \Queue_reg[4][14]  ( .D(n392), .CPN(Clk_r), .Q(\Queue[4][14] ) );
  FDN1QM1P \Queue_reg[3][14]  ( .D(n520), .CPN(Clk_r), .Q(\Queue[3][14] ) );
  FDN1QM1P \Queue_reg[2][14]  ( .D(n488), .CPN(Clk_r), .Q(\Queue[2][14] ) );
  FDN1QM1P \Queue_reg[4][13]  ( .D(n391), .CPN(Clk_r), .Q(\Queue[4][13] ) );
  FDN1QM1P \Queue_reg[3][13]  ( .D(n519), .CPN(Clk_r), .Q(\Queue[3][13] ) );
  FDN1QM1P \Queue_reg[2][13]  ( .D(n487), .CPN(Clk_r), .Q(\Queue[2][13] ) );
  FDN1QM1P \Queue_reg[4][12]  ( .D(n390), .CPN(Clk_r), .Q(\Queue[4][12] ) );
  FDN1QM1P \Queue_reg[3][12]  ( .D(n518), .CPN(Clk_r), .Q(\Queue[3][12] ) );
  FDN1QM1P \Queue_reg[2][12]  ( .D(n486), .CPN(Clk_r), .Q(\Queue[2][12] ) );
  FDN1QM1P \Queue_reg[4][11]  ( .D(n389), .CPN(Clk_r), .Q(\Queue[4][11] ) );
  FDN1QM1P \Queue_reg[3][11]  ( .D(n517), .CPN(Clk_r), .Q(\Queue[3][11] ) );
  FDN1QM1P \Queue_reg[2][11]  ( .D(n485), .CPN(Clk_r), .Q(\Queue[2][11] ) );
  FDN1QM1P \Queue_reg[4][10]  ( .D(n388), .CPN(Clk_r), .Q(\Queue[4][10] ) );
  FDN1QM1P \Queue_reg[3][10]  ( .D(n516), .CPN(Clk_r), .Q(\Queue[3][10] ) );
  FDN1QM1P \Queue_reg[2][10]  ( .D(n484), .CPN(Clk_r), .Q(\Queue[2][10] ) );
  FDN1QM1P \Queue_reg[4][9]  ( .D(n387), .CPN(Clk_r), .Q(\Queue[4][9] ) );
  FDN1QM1P \Queue_reg[3][9]  ( .D(n515), .CPN(Clk_r), .Q(\Queue[3][9] ) );
  FDN1QM1P \Queue_reg[2][9]  ( .D(n483), .CPN(Clk_r), .Q(\Queue[2][9] ) );
  FDN1QM1P \Queue_reg[4][8]  ( .D(n386), .CPN(Clk_r), .Q(\Queue[4][8] ) );
  FDN1QM1P \Queue_reg[3][8]  ( .D(n514), .CPN(Clk_r), .Q(\Queue[3][8] ) );
  FDN1QM1P \Queue_reg[2][8]  ( .D(n482), .CPN(Clk_r), .Q(\Queue[2][8] ) );
  FDN1QM1P \Queue_reg[4][7]  ( .D(n385), .CPN(Clk_r), .Q(\Queue[4][7] ) );
  FDN1QM1P \Queue_reg[3][7]  ( .D(n513), .CPN(Clk_r), .Q(\Queue[3][7] ) );
  FDN1QM1P \Queue_reg[2][7]  ( .D(n481), .CPN(Clk_r), .Q(\Queue[2][7] ) );
  FDN1QM1P \Queue_reg[4][6]  ( .D(n384), .CPN(Clk_r), .Q(\Queue[4][6] ) );
  FDN1QM1P \Queue_reg[3][6]  ( .D(n512), .CPN(Clk_r), .Q(\Queue[3][6] ) );
  FDN1QM1P \Queue_reg[2][6]  ( .D(n480), .CPN(Clk_r), .Q(\Queue[2][6] ) );
  FDN1QM1P \Queue_reg[4][5]  ( .D(n383), .CPN(Clk_r), .Q(\Queue[4][5] ) );
  FDN1QM1P \Queue_reg[3][5]  ( .D(n511), .CPN(Clk_r), .Q(\Queue[3][5] ) );
  FDN1QM1P \Queue_reg[2][5]  ( .D(n479), .CPN(Clk_r), .Q(\Queue[2][5] ) );
  FDN1QM1P \Queue_reg[4][4]  ( .D(n382), .CPN(Clk_r), .Q(\Queue[4][4] ) );
  FDN1QM1P \Queue_reg[3][4]  ( .D(n510), .CPN(Clk_r), .Q(\Queue[3][4] ) );
  FDN1QM1P \Queue_reg[2][4]  ( .D(n478), .CPN(Clk_r), .Q(\Queue[2][4] ) );
  FDN1QM1P \Queue_reg[4][3]  ( .D(n381), .CPN(Clk_r), .Q(\Queue[4][3] ) );
  FDN1QM1P \Queue_reg[3][3]  ( .D(n509), .CPN(Clk_r), .Q(\Queue[3][3] ) );
  FDN1QM1P \Queue_reg[2][3]  ( .D(n477), .CPN(Clk_r), .Q(\Queue[2][3] ) );
  FDN1QM1P \Queue_reg[4][2]  ( .D(n380), .CPN(Clk_r), .Q(\Queue[4][2] ) );
  FDN1QM1P \Queue_reg[3][2]  ( .D(n508), .CPN(Clk_r), .Q(\Queue[3][2] ) );
  FDN1QM1P \Queue_reg[2][2]  ( .D(n476), .CPN(Clk_r), .Q(\Queue[2][2] ) );
  FDN1QM1P \Queue_reg[4][1]  ( .D(n379), .CPN(Clk_r), .Q(\Queue[4][1] ) );
  FDN1QM1P \Queue_reg[3][1]  ( .D(n507), .CPN(Clk_r), .Q(\Queue[3][1] ) );
  FDN1QM1P \Queue_reg[2][1]  ( .D(n475), .CPN(Clk_r), .Q(\Queue[2][1] ) );
  FDN1QM1P \Queue_reg[4][0]  ( .D(n378), .CPN(Clk_r), .Q(\Queue[4][0] ) );
  FDN1QM1P \Queue_reg[3][0]  ( .D(n506), .CPN(Clk_r), .Q(\Queue[3][0] ) );
  FDN1QM1P \Queue_reg[2][0]  ( .D(n474), .CPN(Clk_r), .Q(\Queue[2][0] ) );
  FDN1QM1P \Queue_reg[4][31]  ( .D(n377), .CPN(Clk_r), .Q(\Queue[4][31] ) );
  FDN1QM1P \Queue_reg[3][31]  ( .D(n537), .CPN(Clk_r), .Q(\Queue[3][31] ) );
  FDN1QM1P \Queue_reg[2][31]  ( .D(n505), .CPN(Clk_r), .Q(\Queue[2][31] ) );
  FDN2QM1P Full_reg ( .D(n409), .CPN(Clk_r), .CD(Rst_n), .Q(Full) );
  FDN1QM1P \Queue_reg[1][31]  ( .D(n441), .CPN(Clk_r), .Q(\Queue[1][31] ) );
  FDN1QM1P \Queue_reg[0][31]  ( .D(n473), .CPN(Clk_r), .Q(Packet_Out[31]) );
  FDN1QM1P \Queue_reg[1][30]  ( .D(n440), .CPN(Clk_r), .Q(\Queue[1][30] ) );
  FDN1QM1P \Queue_reg[0][30]  ( .D(n472), .CPN(Clk_r), .Q(Packet_Out[30]) );
  FDN1QM1P \Queue_reg[1][29]  ( .D(n439), .CPN(Clk_r), .Q(\Queue[1][29] ) );
  FDN1QM1P \Queue_reg[0][29]  ( .D(n471), .CPN(Clk_r), .Q(Packet_Out[29]) );
  FDN1QM1P \Queue_reg[1][28]  ( .D(n438), .CPN(Clk_r), .Q(\Queue[1][28] ) );
  FDN1QM1P \Queue_reg[0][28]  ( .D(n470), .CPN(Clk_r), .Q(Packet_Out[28]) );
  FDN1QM1P \Queue_reg[1][27]  ( .D(n437), .CPN(Clk_r), .Q(\Queue[1][27] ) );
  FDN1QM1P \Queue_reg[0][27]  ( .D(n469), .CPN(Clk_r), .Q(Packet_Out[27]) );
  FDN1QM1P \Queue_reg[1][26]  ( .D(n436), .CPN(Clk_r), .Q(\Queue[1][26] ) );
  FDN1QM1P \Queue_reg[0][26]  ( .D(n468), .CPN(Clk_r), .Q(Packet_Out[26]) );
  FDN1QM1P \Queue_reg[1][25]  ( .D(n435), .CPN(Clk_r), .Q(\Queue[1][25] ) );
  FDN1QM1P \Queue_reg[0][25]  ( .D(n467), .CPN(Clk_r), .Q(Packet_Out[25]) );
  FDN1QM1P \Queue_reg[1][24]  ( .D(n434), .CPN(Clk_r), .Q(\Queue[1][24] ) );
  FDN1QM1P \Queue_reg[0][24]  ( .D(n466), .CPN(Clk_r), .Q(Packet_Out[24]) );
  FDN1QM1P \Queue_reg[1][23]  ( .D(n433), .CPN(Clk_r), .Q(\Queue[1][23] ) );
  FDN1QM1P \Queue_reg[0][23]  ( .D(n465), .CPN(Clk_r), .Q(Packet_Out[23]) );
  FDN1QM1P \Queue_reg[1][22]  ( .D(n432), .CPN(Clk_r), .Q(\Queue[1][22] ) );
  FDN1QM1P \Queue_reg[0][22]  ( .D(n464), .CPN(Clk_r), .Q(Packet_Out[22]) );
  FDN1QM1P \Queue_reg[1][21]  ( .D(n431), .CPN(Clk_r), .Q(\Queue[1][21] ) );
  FDN1QM1P \Queue_reg[0][21]  ( .D(n463), .CPN(Clk_r), .Q(Packet_Out[21]) );
  FDN1QM1P \Queue_reg[1][20]  ( .D(n430), .CPN(Clk_r), .Q(\Queue[1][20] ) );
  FDN1QM1P \Queue_reg[0][20]  ( .D(n462), .CPN(Clk_r), .Q(Packet_Out[20]) );
  FDN1QM1P \Queue_reg[1][19]  ( .D(n429), .CPN(Clk_r), .Q(\Queue[1][19] ) );
  FDN1QM1P \Queue_reg[0][19]  ( .D(n461), .CPN(Clk_r), .Q(Packet_Out[19]) );
  FDN1QM1P \Queue_reg[1][18]  ( .D(n428), .CPN(Clk_r), .Q(\Queue[1][18] ) );
  FDN1QM1P \Queue_reg[0][18]  ( .D(n460), .CPN(Clk_r), .Q(Packet_Out[18]) );
  FDN1QM1P \Queue_reg[1][17]  ( .D(n427), .CPN(Clk_r), .Q(\Queue[1][17] ) );
  FDN1QM1P \Queue_reg[0][17]  ( .D(n459), .CPN(Clk_r), .Q(Packet_Out[17]) );
  FDN1QM1P \Queue_reg[1][16]  ( .D(n426), .CPN(Clk_r), .Q(\Queue[1][16] ) );
  FDN1QM1P \Queue_reg[0][16]  ( .D(n458), .CPN(Clk_r), .Q(Packet_Out[16]) );
  FDN1QM1P \Queue_reg[1][15]  ( .D(n425), .CPN(Clk_r), .Q(\Queue[1][15] ) );
  FDN1QM1P \Queue_reg[0][15]  ( .D(n457), .CPN(Clk_r), .Q(Packet_Out[15]) );
  FDN1QM1P \Queue_reg[1][14]  ( .D(n424), .CPN(Clk_r), .Q(\Queue[1][14] ) );
  FDN1QM1P \Queue_reg[0][14]  ( .D(n456), .CPN(Clk_r), .Q(Packet_Out[14]) );
  FDN1QM1P \Queue_reg[1][13]  ( .D(n423), .CPN(Clk_r), .Q(\Queue[1][13] ) );
  FDN1QM1P \Queue_reg[0][13]  ( .D(n455), .CPN(Clk_r), .Q(Packet_Out[13]) );
  FDN1QM1P \Queue_reg[1][12]  ( .D(n422), .CPN(Clk_r), .Q(\Queue[1][12] ) );
  FDN1QM1P \Queue_reg[0][12]  ( .D(n454), .CPN(Clk_r), .Q(Packet_Out[12]) );
  FDN1QM1P \Queue_reg[1][11]  ( .D(n421), .CPN(Clk_r), .Q(\Queue[1][11] ) );
  FDN1QM1P \Queue_reg[0][11]  ( .D(n453), .CPN(Clk_r), .Q(Packet_Out[11]) );
  FDN1QM1P \Queue_reg[1][10]  ( .D(n420), .CPN(Clk_r), .Q(\Queue[1][10] ) );
  FDN1QM1P \Queue_reg[0][10]  ( .D(n452), .CPN(Clk_r), .Q(Packet_Out[10]) );
  FDN1QM1P \Queue_reg[1][9]  ( .D(n419), .CPN(Clk_r), .Q(\Queue[1][9] ) );
  FDN1QM1P \Queue_reg[0][9]  ( .D(n451), .CPN(Clk_r), .Q(Packet_Out[9]) );
  FDN1QM1P \Queue_reg[1][8]  ( .D(n418), .CPN(Clk_r), .Q(\Queue[1][8] ) );
  FDN1QM1P \Queue_reg[0][8]  ( .D(n450), .CPN(Clk_r), .Q(Packet_Out[8]) );
  FDN1QM1P \Queue_reg[1][7]  ( .D(n417), .CPN(Clk_r), .Q(\Queue[1][7] ) );
  FDN1QM1P \Queue_reg[0][7]  ( .D(n449), .CPN(Clk_r), .Q(Packet_Out[7]) );
  FDN1QM1P \Queue_reg[1][6]  ( .D(n416), .CPN(Clk_r), .Q(\Queue[1][6] ) );
  FDN1QM1P \Queue_reg[0][6]  ( .D(n448), .CPN(Clk_r), .Q(Packet_Out[6]) );
  FDN1QM1P \Queue_reg[1][5]  ( .D(n415), .CPN(Clk_r), .Q(\Queue[1][5] ) );
  FDN1QM1P \Queue_reg[0][5]  ( .D(n447), .CPN(Clk_r), .Q(Packet_Out[5]) );
  FDN1QM1P \Queue_reg[1][4]  ( .D(n414), .CPN(Clk_r), .Q(\Queue[1][4] ) );
  FDN1QM1P \Queue_reg[0][4]  ( .D(n446), .CPN(Clk_r), .Q(Packet_Out[4]) );
  FDN1QM1P \Queue_reg[1][3]  ( .D(n413), .CPN(Clk_r), .Q(\Queue[1][3] ) );
  FDN1QM1P \Queue_reg[0][3]  ( .D(n445), .CPN(Clk_r), .Q(Packet_Out[3]) );
  FDN1QM1P \Queue_reg[1][2]  ( .D(n412), .CPN(Clk_r), .Q(\Queue[1][2] ) );
  FDN1QM1P \Queue_reg[0][2]  ( .D(n444), .CPN(Clk_r), .Q(Packet_Out[2]) );
  FDN1QM1P \Queue_reg[1][1]  ( .D(n411), .CPN(Clk_r), .Q(\Queue[1][1] ) );
  FDN1QM1P \Queue_reg[0][1]  ( .D(n443), .CPN(Clk_r), .Q(Packet_Out[1]) );
  FDN1QM1P \Queue_reg[1][0]  ( .D(n410), .CPN(Clk_r), .Q(\Queue[1][0] ) );
  FDN1QM1P \Queue_reg[0][0]  ( .D(n442), .CPN(Clk_r), .Q(Packet_Out[0]) );
  FDN2QM1P Empty_reg ( .D(n539), .CPN(Clk_r), .CD(Rst_n), .Q(n538) );
  BUFM3P U3 ( .A(n94), .Z(n9) );
  OAI211M4P U4 ( .A(n97), .B(n134), .C(Write_Ack), .D(n22), .Z(n3) );
  AOI21M3P U5 ( .A(Write_Ack), .B(n139), .C(n138), .Z(n202) );
  N1M1P U6 ( .A(Read_Ack), .Z(n134) );
  N1M1P U7 ( .A(Write_Ack), .Z(n96) );
  AOI21M3P U8 ( .A(Write_Ack), .B(n97), .C(n138), .Z(n55) );
  OAI211M4P U9 ( .A(n137), .B(n136), .C(Rst_n), .D(n135), .Z(n203) );
  AOI21M3P U10 ( .A(Write_Ack), .B(n373), .C(n138), .Z(n92) );
  OAI211M4P U11 ( .A(n97), .B(n136), .C(Rst_n), .D(n135), .Z(n130) );
  NR2I1M8P U12 ( .A(n58), .B(n19), .Z(n18) );
  AOI21M3P U13 ( .A(Write_Ack), .B(n137), .C(n138), .Z(n129) );
  ND2M1P U14 ( .A(n16), .B(Rst_n), .Z(n58) );
  NR2M2P U15 ( .A(Read_Ack), .B(n96), .Z(n16) );
  NR3M1P U16 ( .A(Count[2]), .B(n21), .C(n20), .Z(n137) );
  NR3M1P U17 ( .A(Count[0]), .B(Count[1]), .C(n17), .Z(n139) );
  NR3M1P U18 ( .A(n21), .B(Count[2]), .C(Count[1]), .Z(n373) );
  NR3M1P U19 ( .A(Count[0]), .B(Count[2]), .C(n20), .Z(n97) );
  N1M1P U20 ( .A(Count[1]), .Z(n20) );
  N1M1P U21 ( .A(Count[0]), .Z(n21) );
  N1M1P U22 ( .A(Count[2]), .Z(n17) );
  ND2M2P U23 ( .A(Read_Ack), .B(Rst_n), .Z(n138) );
  OAI211M4P U24 ( .A(n139), .B(n134), .C(Write_Ack), .D(n133), .Z(n205) );
  BUFM2P U25 ( .A(n91), .Z(n7) );
  BUFM2P U26 ( .A(n91), .Z(n8) );
  N1M2P U27 ( .A(n59), .Z(n91) );
  BUFM2P U28 ( .A(n94), .Z(n10) );
  OAI211M1P U29 ( .A(n373), .B(n134), .C(Write_Ack), .D(n59), .Z(n94) );
  BUFM2P U30 ( .A(n54), .Z(n5) );
  BUFM2P U31 ( .A(n54), .Z(n4) );
  BUFM2P U32 ( .A(n54), .Z(n6) );
  N1M2P U33 ( .A(n16), .Z(n136) );
  OAI211M4P U34 ( .A(n137), .B(n134), .C(Write_Ack), .D(n95), .Z(n132) );
  AOI22M1P U35 ( .A(Count[0]), .B(n136), .C(n15), .D(n21), .Z(n12) );
  NR2M1P U36 ( .A(n134), .B(Write_Ack), .Z(n208) );
  NR2M1P U37 ( .A(n16), .B(n208), .Z(n207) );
  AOI22CDNM1P U38 ( .A(n207), .B(n21), .C(n207), .D(n21), .Z(n374) );
  N1M1P U39 ( .A(n208), .Z(n15) );
  AOI22CDNM1P U40 ( .A(Count[1]), .B(n12), .C(n12), .D(Count[1]), .Z(n375) );
  ND3M1P U41 ( .A(n21), .B(n17), .C(n20), .Z(n57) );
  ND2M1P U42 ( .A(Count[1]), .B(Read_Ack), .Z(n11) );
  OAI211M1P U43 ( .A(Count[1]), .B(n136), .C(n12), .D(n11), .Z(n13) );
  AOI22M1P U44 ( .A(n16), .B(n137), .C(Count[2]), .D(n13), .Z(n14) );
  OAI21M1P U45 ( .A(n57), .B(n15), .C(n14), .Z(n376) );
  N1M1P U46 ( .A(n139), .Z(n19) );
  N1M1P U47 ( .A(Packet_In[31]), .Z(n206) );
  AOI22CDNM1P U48 ( .A(n18), .B(n206), .C(\Queue[4][31] ), .D(n18), .Z(n377)
         );
  N1M1P U49 ( .A(Packet_In[0]), .Z(n141) );
  AOI22CDNM1P U50 ( .A(n18), .B(n141), .C(\Queue[4][0] ), .D(n18), .Z(n378) );
  N1M1P U51 ( .A(Packet_In[1]), .Z(n143) );
  AOI22CDNM1P U52 ( .A(n18), .B(n143), .C(\Queue[4][1] ), .D(n18), .Z(n379) );
  N1M1P U53 ( .A(Packet_In[2]), .Z(n145) );
  AOI22CDNM1P U54 ( .A(n18), .B(n145), .C(\Queue[4][2] ), .D(n18), .Z(n380) );
  N1M1P U55 ( .A(Packet_In[3]), .Z(n147) );
  AOI22CDNM1P U56 ( .A(n18), .B(n147), .C(\Queue[4][3] ), .D(n18), .Z(n381) );
  N1M1P U57 ( .A(Packet_In[4]), .Z(n149) );
  AOI22CDNM1P U58 ( .A(n18), .B(n149), .C(\Queue[4][4] ), .D(n18), .Z(n382) );
  N1M1P U59 ( .A(Packet_In[5]), .Z(n151) );
  AOI22CDNM1P U60 ( .A(n18), .B(n151), .C(\Queue[4][5] ), .D(n18), .Z(n383) );
  N1M1P U61 ( .A(Packet_In[6]), .Z(n153) );
  AOI22CDNM1P U62 ( .A(n18), .B(n153), .C(\Queue[4][6] ), .D(n18), .Z(n384) );
  N1M1P U63 ( .A(Packet_In[7]), .Z(n155) );
  AOI22CDNM1P U64 ( .A(n18), .B(n155), .C(\Queue[4][7] ), .D(n18), .Z(n385) );
  N1M1P U65 ( .A(Packet_In[8]), .Z(n157) );
  AOI22CDNM1P U66 ( .A(n18), .B(n157), .C(\Queue[4][8] ), .D(n18), .Z(n386) );
  N1M1P U67 ( .A(Packet_In[9]), .Z(n159) );
  AOI22CDNM1P U68 ( .A(n18), .B(n159), .C(\Queue[4][9] ), .D(n18), .Z(n387) );
  N1M1P U69 ( .A(Packet_In[10]), .Z(n161) );
  AOI22CDNM1P U70 ( .A(n18), .B(n161), .C(\Queue[4][10] ), .D(n18), .Z(n388)
         );
  N1M1P U71 ( .A(Packet_In[11]), .Z(n163) );
  AOI22CDNM1P U72 ( .A(n18), .B(n163), .C(\Queue[4][11] ), .D(n18), .Z(n389)
         );
  N1M1P U73 ( .A(Packet_In[12]), .Z(n165) );
  AOI22CDNM1P U74 ( .A(n18), .B(n165), .C(\Queue[4][12] ), .D(n18), .Z(n390)
         );
  N1M1P U75 ( .A(Packet_In[13]), .Z(n167) );
  AOI22CDNM1P U76 ( .A(n18), .B(n167), .C(\Queue[4][13] ), .D(n18), .Z(n391)
         );
  N1M1P U77 ( .A(Packet_In[14]), .Z(n169) );
  AOI22CDNM1P U78 ( .A(n18), .B(n169), .C(\Queue[4][14] ), .D(n18), .Z(n392)
         );
  N1M1P U79 ( .A(Packet_In[15]), .Z(n171) );
  AOI22CDNM1P U80 ( .A(n18), .B(n171), .C(\Queue[4][15] ), .D(n18), .Z(n393)
         );
  N1M1P U81 ( .A(Packet_In[16]), .Z(n173) );
  AOI22CDNM1P U82 ( .A(n18), .B(n173), .C(\Queue[4][16] ), .D(n18), .Z(n394)
         );
  N1M1P U83 ( .A(Packet_In[17]), .Z(n175) );
  AOI22CDNM1P U84 ( .A(n18), .B(n175), .C(\Queue[4][17] ), .D(n18), .Z(n395)
         );
  N1M1P U85 ( .A(Packet_In[18]), .Z(n177) );
  AOI22CDNM1P U86 ( .A(n18), .B(n177), .C(\Queue[4][18] ), .D(n18), .Z(n396)
         );
  N1M1P U87 ( .A(Packet_In[19]), .Z(n179) );
  AOI22CDNM1P U88 ( .A(n18), .B(n179), .C(\Queue[4][19] ), .D(n18), .Z(n397)
         );
  N1M1P U89 ( .A(Packet_In[20]), .Z(n181) );
  AOI22CDNM1P U90 ( .A(n18), .B(n181), .C(\Queue[4][20] ), .D(n18), .Z(n398)
         );
  N1M1P U91 ( .A(Packet_In[21]), .Z(n183) );
  AOI22CDNM1P U92 ( .A(n18), .B(n183), .C(\Queue[4][21] ), .D(n18), .Z(n399)
         );
  N1M1P U93 ( .A(Packet_In[22]), .Z(n185) );
  AOI22CDNM1P U94 ( .A(n18), .B(n185), .C(\Queue[4][22] ), .D(n18), .Z(n400)
         );
  N1M1P U95 ( .A(Packet_In[23]), .Z(n187) );
  AOI22CDNM1P U96 ( .A(n18), .B(n187), .C(\Queue[4][23] ), .D(n18), .Z(n401)
         );
  N1M1P U97 ( .A(Packet_In[24]), .Z(n189) );
  AOI22CDNM1P U98 ( .A(n18), .B(n189), .C(\Queue[4][24] ), .D(n18), .Z(n402)
         );
  N1M1P U99 ( .A(Packet_In[25]), .Z(n191) );
  AOI22CDNM1P U100 ( .A(n18), .B(n191), .C(\Queue[4][25] ), .D(n18), .Z(n403)
         );
  N1M1P U101 ( .A(Packet_In[26]), .Z(n193) );
  AOI22CDNM1P U102 ( .A(n18), .B(n193), .C(\Queue[4][26] ), .D(n18), .Z(n404)
         );
  N1M1P U103 ( .A(Packet_In[27]), .Z(n195) );
  AOI22CDNM1P U104 ( .A(n18), .B(n195), .C(\Queue[4][27] ), .D(n18), .Z(n405)
         );
  N1M1P U105 ( .A(Packet_In[28]), .Z(n197) );
  AOI22CDNM1P U106 ( .A(n18), .B(n197), .C(\Queue[4][28] ), .D(n18), .Z(n406)
         );
  N1M1P U107 ( .A(Packet_In[29]), .Z(n199) );
  AOI22CDNM1P U108 ( .A(n18), .B(n199), .C(\Queue[4][29] ), .D(n18), .Z(n407)
         );
  N1M1P U109 ( .A(Packet_In[30]), .Z(n201) );
  AOI22CDNM1P U110 ( .A(n18), .B(n201), .C(\Queue[4][30] ), .D(n18), .Z(n408)
         );
  OAI22CDNM1P U111 ( .A(n136), .B(n19), .C(n207), .D(Full), .Z(n409) );
  OA21M1P U112 ( .A(n136), .B(n373), .C(Rst_n), .Z(n22) );
  OAI21M1P U113 ( .A(Write_Ack), .B(Read_Ack), .C(n22), .Z(n54) );
  AOI22M1P U114 ( .A(\Queue[2][0] ), .B(n55), .C(\Queue[1][0] ), .D(n4), .Z(
        n23) );
  OAI21M1P U115 ( .A(n141), .B(n3), .C(n23), .Z(n410) );
  AOI22M1P U116 ( .A(n55), .B(\Queue[2][1] ), .C(\Queue[1][1] ), .D(n4), .Z(
        n24) );
  OAI21M1P U117 ( .A(n3), .B(n143), .C(n24), .Z(n411) );
  AOI22M1P U118 ( .A(n55), .B(\Queue[2][2] ), .C(\Queue[1][2] ), .D(n4), .Z(
        n25) );
  OAI21M1P U119 ( .A(n3), .B(n145), .C(n25), .Z(n412) );
  AOI22M1P U120 ( .A(n55), .B(\Queue[2][3] ), .C(\Queue[1][3] ), .D(n4), .Z(
        n26) );
  OAI21M1P U121 ( .A(n3), .B(n147), .C(n26), .Z(n413) );
  AOI22M1P U122 ( .A(n55), .B(\Queue[2][4] ), .C(\Queue[1][4] ), .D(n4), .Z(
        n27) );
  OAI21M1P U123 ( .A(n3), .B(n149), .C(n27), .Z(n414) );
  AOI22M1P U124 ( .A(n55), .B(\Queue[2][5] ), .C(\Queue[1][5] ), .D(n4), .Z(
        n28) );
  OAI21M1P U125 ( .A(n3), .B(n151), .C(n28), .Z(n415) );
  AOI22M1P U126 ( .A(n55), .B(\Queue[2][6] ), .C(\Queue[1][6] ), .D(n4), .Z(
        n29) );
  OAI21M1P U127 ( .A(n3), .B(n153), .C(n29), .Z(n416) );
  AOI22M1P U128 ( .A(n55), .B(\Queue[2][7] ), .C(\Queue[1][7] ), .D(n4), .Z(
        n30) );
  OAI21M1P U129 ( .A(n3), .B(n155), .C(n30), .Z(n417) );
  AOI22M1P U130 ( .A(n55), .B(\Queue[2][8] ), .C(\Queue[1][8] ), .D(n4), .Z(
        n31) );
  OAI21M1P U131 ( .A(n3), .B(n157), .C(n31), .Z(n418) );
  AOI22M1P U132 ( .A(n55), .B(\Queue[2][9] ), .C(\Queue[1][9] ), .D(n5), .Z(
        n32) );
  OAI21M1P U133 ( .A(n3), .B(n159), .C(n32), .Z(n419) );
  AOI22M1P U134 ( .A(n55), .B(\Queue[2][10] ), .C(\Queue[1][10] ), .D(n5), .Z(
        n33) );
  OAI21M1P U135 ( .A(n3), .B(n161), .C(n33), .Z(n420) );
  AOI22M1P U136 ( .A(n55), .B(\Queue[2][11] ), .C(\Queue[1][11] ), .D(n5), .Z(
        n34) );
  OAI21M1P U137 ( .A(n3), .B(n163), .C(n34), .Z(n421) );
  AOI22M1P U138 ( .A(n55), .B(\Queue[2][12] ), .C(\Queue[1][12] ), .D(n5), .Z(
        n35) );
  OAI21M1P U139 ( .A(n3), .B(n165), .C(n35), .Z(n422) );
  AOI22M1P U140 ( .A(n55), .B(\Queue[2][13] ), .C(\Queue[1][13] ), .D(n5), .Z(
        n36) );
  OAI21M1P U141 ( .A(n3), .B(n167), .C(n36), .Z(n423) );
  AOI22M1P U142 ( .A(n55), .B(\Queue[2][14] ), .C(\Queue[1][14] ), .D(n5), .Z(
        n37) );
  OAI21M1P U143 ( .A(n3), .B(n169), .C(n37), .Z(n424) );
  AOI22M1P U144 ( .A(n55), .B(\Queue[2][15] ), .C(\Queue[1][15] ), .D(n5), .Z(
        n38) );
  OAI21M1P U145 ( .A(n3), .B(n171), .C(n38), .Z(n425) );
  AOI22M1P U146 ( .A(n55), .B(\Queue[2][16] ), .C(\Queue[1][16] ), .D(n5), .Z(
        n39) );
  OAI21M1P U147 ( .A(n3), .B(n173), .C(n39), .Z(n426) );
  AOI22M1P U148 ( .A(n55), .B(\Queue[2][17] ), .C(\Queue[1][17] ), .D(n5), .Z(
        n40) );
  OAI21M1P U149 ( .A(n3), .B(n175), .C(n40), .Z(n427) );
  AOI22M1P U150 ( .A(n55), .B(\Queue[2][18] ), .C(\Queue[1][18] ), .D(n6), .Z(
        n41) );
  OAI21M1P U151 ( .A(n3), .B(n177), .C(n41), .Z(n428) );
  AOI22M1P U152 ( .A(n55), .B(\Queue[2][19] ), .C(\Queue[1][19] ), .D(n6), .Z(
        n42) );
  OAI21M1P U153 ( .A(n3), .B(n179), .C(n42), .Z(n429) );
  AOI22M1P U154 ( .A(n55), .B(\Queue[2][20] ), .C(\Queue[1][20] ), .D(n6), .Z(
        n43) );
  OAI21M1P U155 ( .A(n3), .B(n181), .C(n43), .Z(n430) );
  AOI22M1P U156 ( .A(n55), .B(\Queue[2][21] ), .C(\Queue[1][21] ), .D(n6), .Z(
        n44) );
  OAI21M1P U157 ( .A(n3), .B(n183), .C(n44), .Z(n431) );
  AOI22M1P U158 ( .A(n55), .B(\Queue[2][22] ), .C(\Queue[1][22] ), .D(n6), .Z(
        n45) );
  OAI21M1P U159 ( .A(n3), .B(n185), .C(n45), .Z(n432) );
  AOI22M1P U160 ( .A(n55), .B(\Queue[2][23] ), .C(\Queue[1][23] ), .D(n6), .Z(
        n46) );
  OAI21M1P U161 ( .A(n3), .B(n187), .C(n46), .Z(n433) );
  AOI22M1P U162 ( .A(n55), .B(\Queue[2][24] ), .C(\Queue[1][24] ), .D(n6), .Z(
        n47) );
  OAI21M1P U163 ( .A(n3), .B(n189), .C(n47), .Z(n434) );
  AOI22M1P U164 ( .A(n55), .B(\Queue[2][25] ), .C(\Queue[1][25] ), .D(n6), .Z(
        n48) );
  OAI21M1P U165 ( .A(n3), .B(n191), .C(n48), .Z(n435) );
  AOI22M1P U166 ( .A(n55), .B(\Queue[2][26] ), .C(\Queue[1][26] ), .D(n6), .Z(
        n49) );
  OAI21M1P U167 ( .A(n3), .B(n193), .C(n49), .Z(n436) );
  AOI22M1P U168 ( .A(n55), .B(\Queue[2][27] ), .C(\Queue[1][27] ), .D(n6), .Z(
        n50) );
  OAI21M1P U169 ( .A(n3), .B(n195), .C(n50), .Z(n437) );
  AOI22M1P U170 ( .A(n55), .B(\Queue[2][28] ), .C(\Queue[1][28] ), .D(n4), .Z(
        n51) );
  OAI21M1P U171 ( .A(n3), .B(n197), .C(n51), .Z(n438) );
  AOI22M1P U172 ( .A(n55), .B(\Queue[2][29] ), .C(\Queue[1][29] ), .D(n5), .Z(
        n52) );
  OAI21M1P U173 ( .A(n3), .B(n199), .C(n52), .Z(n439) );
  AOI22M1P U174 ( .A(n55), .B(\Queue[2][30] ), .C(\Queue[1][30] ), .D(n6), .Z(
        n53) );
  OAI21M1P U175 ( .A(n3), .B(n201), .C(n53), .Z(n440) );
  AOI22M1P U176 ( .A(n55), .B(\Queue[2][31] ), .C(\Queue[1][31] ), .D(n4), .Z(
        n56) );
  OAI21M1P U177 ( .A(n3), .B(n206), .C(n56), .Z(n441) );
  OAI21M1P U178 ( .A(n58), .B(n57), .C(n138), .Z(n59) );
  AOI22M1P U179 ( .A(\Queue[1][0] ), .B(n92), .C(n91), .D(Packet_Out[0]), .Z(
        n60) );
  OAI21M1P U180 ( .A(n141), .B(n9), .C(n60), .Z(n442) );
  AOI22M1P U181 ( .A(\Queue[1][1] ), .B(n92), .C(n91), .D(Packet_Out[1]), .Z(
        n61) );
  OAI21M1P U182 ( .A(n143), .B(n9), .C(n61), .Z(n443) );
  AOI22M1P U183 ( .A(\Queue[1][2] ), .B(n92), .C(n91), .D(Packet_Out[2]), .Z(
        n62) );
  OAI21M1P U184 ( .A(n145), .B(n9), .C(n62), .Z(n444) );
  AOI22M1P U185 ( .A(\Queue[1][3] ), .B(n92), .C(n91), .D(Packet_Out[3]), .Z(
        n63) );
  OAI21M1P U186 ( .A(n147), .B(n9), .C(n63), .Z(n445) );
  AOI22M1P U187 ( .A(\Queue[1][4] ), .B(n92), .C(n91), .D(Packet_Out[4]), .Z(
        n64) );
  OAI21M1P U188 ( .A(n149), .B(n9), .C(n64), .Z(n446) );
  AOI22M1P U189 ( .A(\Queue[1][5] ), .B(n92), .C(n91), .D(Packet_Out[5]), .Z(
        n65) );
  OAI21M1P U190 ( .A(n151), .B(n9), .C(n65), .Z(n447) );
  AOI22M1P U191 ( .A(\Queue[1][6] ), .B(n92), .C(n91), .D(Packet_Out[6]), .Z(
        n66) );
  OAI21M1P U192 ( .A(n153), .B(n9), .C(n66), .Z(n448) );
  AOI22M1P U193 ( .A(\Queue[1][7] ), .B(n92), .C(n91), .D(Packet_Out[7]), .Z(
        n67) );
  OAI21M1P U194 ( .A(n155), .B(n9), .C(n67), .Z(n449) );
  AOI22M1P U195 ( .A(\Queue[1][8] ), .B(n92), .C(n91), .D(Packet_Out[8]), .Z(
        n68) );
  OAI21M1P U196 ( .A(n157), .B(n9), .C(n68), .Z(n450) );
  AOI22M1P U197 ( .A(\Queue[1][9] ), .B(n92), .C(n91), .D(Packet_Out[9]), .Z(
        n69) );
  OAI21M1P U198 ( .A(n159), .B(n9), .C(n69), .Z(n451) );
  AOI22M1P U199 ( .A(\Queue[1][10] ), .B(n92), .C(n7), .D(Packet_Out[10]), .Z(
        n70) );
  OAI21M1P U200 ( .A(n161), .B(n9), .C(n70), .Z(n452) );
  AOI22M1P U201 ( .A(\Queue[1][11] ), .B(n92), .C(n7), .D(Packet_Out[11]), .Z(
        n71) );
  OAI21M1P U202 ( .A(n163), .B(n9), .C(n71), .Z(n453) );
  AOI22M1P U203 ( .A(\Queue[1][12] ), .B(n92), .C(n7), .D(Packet_Out[12]), .Z(
        n72) );
  OAI21M1P U204 ( .A(n165), .B(n9), .C(n72), .Z(n454) );
  AOI22M1P U205 ( .A(\Queue[1][13] ), .B(n92), .C(n7), .D(Packet_Out[13]), .Z(
        n73) );
  OAI21M1P U206 ( .A(n167), .B(n9), .C(n73), .Z(n455) );
  AOI22M1P U207 ( .A(\Queue[1][14] ), .B(n92), .C(n7), .D(Packet_Out[14]), .Z(
        n74) );
  OAI21M1P U208 ( .A(n169), .B(n9), .C(n74), .Z(n456) );
  AOI22M1P U209 ( .A(\Queue[1][15] ), .B(n92), .C(n7), .D(Packet_Out[15]), .Z(
        n75) );
  OAI21M1P U210 ( .A(n171), .B(n9), .C(n75), .Z(n457) );
  AOI22M1P U211 ( .A(\Queue[1][16] ), .B(n92), .C(n7), .D(Packet_Out[16]), .Z(
        n76) );
  OAI21M1P U212 ( .A(n173), .B(n9), .C(n76), .Z(n458) );
  AOI22M1P U213 ( .A(\Queue[1][17] ), .B(n92), .C(n7), .D(Packet_Out[17]), .Z(
        n77) );
  OAI21M1P U214 ( .A(n175), .B(n9), .C(n77), .Z(n459) );
  AOI22M1P U215 ( .A(\Queue[1][18] ), .B(n92), .C(n7), .D(Packet_Out[18]), .Z(
        n78) );
  OAI21M1P U216 ( .A(n177), .B(n9), .C(n78), .Z(n460) );
  AOI22M1P U217 ( .A(\Queue[1][19] ), .B(n92), .C(n7), .D(Packet_Out[19]), .Z(
        n79) );
  OAI21M1P U218 ( .A(n179), .B(n9), .C(n79), .Z(n461) );
  AOI22M1P U219 ( .A(\Queue[1][20] ), .B(n92), .C(n8), .D(Packet_Out[20]), .Z(
        n80) );
  OAI21M1P U220 ( .A(n181), .B(n10), .C(n80), .Z(n462) );
  AOI22M1P U221 ( .A(\Queue[1][21] ), .B(n92), .C(n8), .D(Packet_Out[21]), .Z(
        n81) );
  OAI21M1P U222 ( .A(n183), .B(n10), .C(n81), .Z(n463) );
  AOI22M1P U223 ( .A(\Queue[1][22] ), .B(n92), .C(n8), .D(Packet_Out[22]), .Z(
        n82) );
  OAI21M1P U224 ( .A(n185), .B(n10), .C(n82), .Z(n464) );
  AOI22M1P U225 ( .A(\Queue[1][23] ), .B(n92), .C(n8), .D(Packet_Out[23]), .Z(
        n83) );
  OAI21M1P U226 ( .A(n187), .B(n10), .C(n83), .Z(n465) );
  AOI22M1P U227 ( .A(\Queue[1][24] ), .B(n92), .C(n8), .D(Packet_Out[24]), .Z(
        n84) );
  OAI21M1P U228 ( .A(n189), .B(n10), .C(n84), .Z(n466) );
  AOI22M1P U229 ( .A(\Queue[1][25] ), .B(n92), .C(n8), .D(Packet_Out[25]), .Z(
        n85) );
  OAI21M1P U230 ( .A(n191), .B(n10), .C(n85), .Z(n467) );
  AOI22M1P U231 ( .A(\Queue[1][26] ), .B(n92), .C(n8), .D(Packet_Out[26]), .Z(
        n86) );
  OAI21M1P U232 ( .A(n193), .B(n10), .C(n86), .Z(n468) );
  AOI22M1P U233 ( .A(\Queue[1][27] ), .B(n92), .C(n8), .D(Packet_Out[27]), .Z(
        n87) );
  OAI21M1P U234 ( .A(n195), .B(n10), .C(n87), .Z(n469) );
  AOI22M1P U235 ( .A(\Queue[1][28] ), .B(n92), .C(n8), .D(Packet_Out[28]), .Z(
        n88) );
  OAI21M1P U236 ( .A(n197), .B(n10), .C(n88), .Z(n470) );
  AOI22M1P U237 ( .A(\Queue[1][29] ), .B(n92), .C(n8), .D(Packet_Out[29]), .Z(
        n89) );
  OAI21M1P U238 ( .A(n199), .B(n10), .C(n89), .Z(n471) );
  AOI22M1P U239 ( .A(\Queue[1][30] ), .B(n92), .C(n7), .D(Packet_Out[30]), .Z(
        n90) );
  OAI21M1P U240 ( .A(n201), .B(n9), .C(n90), .Z(n472) );
  AOI22M1P U241 ( .A(\Queue[1][31] ), .B(n92), .C(n8), .D(Packet_Out[31]), .Z(
        n93) );
  OAI21M1P U242 ( .A(n206), .B(n10), .C(n93), .Z(n473) );
  OA21M1P U243 ( .A(n136), .B(n97), .C(Rst_n), .Z(n95) );
  ND2M1P U244 ( .A(n96), .B(n134), .Z(n135) );
  AOI22M1P U245 ( .A(\Queue[2][0] ), .B(n130), .C(\Queue[3][0] ), .D(n129), 
        .Z(n98) );
  OAI21M1P U246 ( .A(n141), .B(n132), .C(n98), .Z(n474) );
  AOI22M1P U247 ( .A(\Queue[2][1] ), .B(n130), .C(n129), .D(\Queue[3][1] ), 
        .Z(n99) );
  OAI21M1P U248 ( .A(n143), .B(n132), .C(n99), .Z(n475) );
  AOI22M1P U249 ( .A(\Queue[2][2] ), .B(n130), .C(n129), .D(\Queue[3][2] ), 
        .Z(n100) );
  OAI21M1P U250 ( .A(n145), .B(n132), .C(n100), .Z(n476) );
  AOI22M1P U251 ( .A(\Queue[2][3] ), .B(n130), .C(n129), .D(\Queue[3][3] ), 
        .Z(n101) );
  OAI21M1P U252 ( .A(n147), .B(n132), .C(n101), .Z(n477) );
  AOI22M1P U253 ( .A(\Queue[2][4] ), .B(n130), .C(n129), .D(\Queue[3][4] ), 
        .Z(n102) );
  OAI21M1P U254 ( .A(n149), .B(n132), .C(n102), .Z(n478) );
  AOI22M1P U255 ( .A(\Queue[2][5] ), .B(n130), .C(n129), .D(\Queue[3][5] ), 
        .Z(n103) );
  OAI21M1P U256 ( .A(n151), .B(n132), .C(n103), .Z(n479) );
  AOI22M1P U257 ( .A(\Queue[2][6] ), .B(n130), .C(n129), .D(\Queue[3][6] ), 
        .Z(n104) );
  OAI21M1P U258 ( .A(n153), .B(n132), .C(n104), .Z(n480) );
  AOI22M1P U259 ( .A(\Queue[2][7] ), .B(n130), .C(n129), .D(\Queue[3][7] ), 
        .Z(n105) );
  OAI21M1P U260 ( .A(n155), .B(n132), .C(n105), .Z(n481) );
  AOI22M1P U261 ( .A(\Queue[2][8] ), .B(n130), .C(n129), .D(\Queue[3][8] ), 
        .Z(n106) );
  OAI21M1P U262 ( .A(n157), .B(n132), .C(n106), .Z(n482) );
  AOI22M1P U263 ( .A(\Queue[2][9] ), .B(n130), .C(n129), .D(\Queue[3][9] ), 
        .Z(n107) );
  OAI21M1P U264 ( .A(n159), .B(n132), .C(n107), .Z(n483) );
  AOI22M1P U265 ( .A(\Queue[2][10] ), .B(n130), .C(n129), .D(\Queue[3][10] ), 
        .Z(n108) );
  OAI21M1P U266 ( .A(n161), .B(n132), .C(n108), .Z(n484) );
  AOI22M1P U267 ( .A(\Queue[2][11] ), .B(n130), .C(n129), .D(\Queue[3][11] ), 
        .Z(n109) );
  OAI21M1P U268 ( .A(n163), .B(n132), .C(n109), .Z(n485) );
  AOI22M1P U269 ( .A(\Queue[2][12] ), .B(n130), .C(n129), .D(\Queue[3][12] ), 
        .Z(n110) );
  OAI21M1P U270 ( .A(n165), .B(n132), .C(n110), .Z(n486) );
  AOI22M1P U271 ( .A(\Queue[2][13] ), .B(n130), .C(n129), .D(\Queue[3][13] ), 
        .Z(n111) );
  OAI21M1P U272 ( .A(n167), .B(n132), .C(n111), .Z(n487) );
  AOI22M1P U273 ( .A(\Queue[2][14] ), .B(n130), .C(n129), .D(\Queue[3][14] ), 
        .Z(n112) );
  OAI21M1P U274 ( .A(n169), .B(n132), .C(n112), .Z(n488) );
  AOI22M1P U275 ( .A(\Queue[2][15] ), .B(n130), .C(n129), .D(\Queue[3][15] ), 
        .Z(n113) );
  OAI21M1P U276 ( .A(n171), .B(n132), .C(n113), .Z(n489) );
  AOI22M1P U277 ( .A(\Queue[2][16] ), .B(n130), .C(n129), .D(\Queue[3][16] ), 
        .Z(n114) );
  OAI21M1P U278 ( .A(n173), .B(n132), .C(n114), .Z(n490) );
  AOI22M1P U279 ( .A(\Queue[2][17] ), .B(n130), .C(n129), .D(\Queue[3][17] ), 
        .Z(n115) );
  OAI21M1P U280 ( .A(n175), .B(n132), .C(n115), .Z(n491) );
  AOI22M1P U281 ( .A(\Queue[2][18] ), .B(n130), .C(n129), .D(\Queue[3][18] ), 
        .Z(n116) );
  OAI21M1P U282 ( .A(n177), .B(n132), .C(n116), .Z(n492) );
  AOI22M1P U283 ( .A(\Queue[2][19] ), .B(n130), .C(n129), .D(\Queue[3][19] ), 
        .Z(n117) );
  OAI21M1P U284 ( .A(n179), .B(n132), .C(n117), .Z(n493) );
  AOI22M1P U285 ( .A(\Queue[2][20] ), .B(n130), .C(n129), .D(\Queue[3][20] ), 
        .Z(n118) );
  OAI21M1P U286 ( .A(n181), .B(n132), .C(n118), .Z(n494) );
  AOI22M1P U287 ( .A(\Queue[2][21] ), .B(n130), .C(n129), .D(\Queue[3][21] ), 
        .Z(n119) );
  OAI21M1P U288 ( .A(n183), .B(n132), .C(n119), .Z(n495) );
  AOI22M1P U289 ( .A(\Queue[2][22] ), .B(n130), .C(n129), .D(\Queue[3][22] ), 
        .Z(n120) );
  OAI21M1P U290 ( .A(n185), .B(n132), .C(n120), .Z(n496) );
  AOI22M1P U291 ( .A(\Queue[2][23] ), .B(n130), .C(n129), .D(\Queue[3][23] ), 
        .Z(n121) );
  OAI21M1P U292 ( .A(n187), .B(n132), .C(n121), .Z(n497) );
  AOI22M1P U293 ( .A(\Queue[2][24] ), .B(n130), .C(n129), .D(\Queue[3][24] ), 
        .Z(n122) );
  OAI21M1P U294 ( .A(n189), .B(n132), .C(n122), .Z(n498) );
  AOI22M1P U295 ( .A(\Queue[2][25] ), .B(n130), .C(n129), .D(\Queue[3][25] ), 
        .Z(n123) );
  OAI21M1P U296 ( .A(n191), .B(n132), .C(n123), .Z(n499) );
  AOI22M1P U297 ( .A(\Queue[2][26] ), .B(n130), .C(n129), .D(\Queue[3][26] ), 
        .Z(n124) );
  OAI21M1P U298 ( .A(n193), .B(n132), .C(n124), .Z(n500) );
  AOI22M1P U299 ( .A(\Queue[2][27] ), .B(n130), .C(n129), .D(\Queue[3][27] ), 
        .Z(n125) );
  OAI21M1P U300 ( .A(n195), .B(n132), .C(n125), .Z(n501) );
  AOI22M1P U301 ( .A(\Queue[2][28] ), .B(n130), .C(n129), .D(\Queue[3][28] ), 
        .Z(n126) );
  OAI21M1P U302 ( .A(n197), .B(n132), .C(n126), .Z(n502) );
  AOI22M1P U303 ( .A(\Queue[2][29] ), .B(n130), .C(n129), .D(\Queue[3][29] ), 
        .Z(n127) );
  OAI21M1P U304 ( .A(n199), .B(n132), .C(n127), .Z(n503) );
  AOI22M1P U305 ( .A(\Queue[2][30] ), .B(n130), .C(n129), .D(\Queue[3][30] ), 
        .Z(n128) );
  OAI21M1P U306 ( .A(n201), .B(n132), .C(n128), .Z(n504) );
  AOI22M1P U307 ( .A(\Queue[2][31] ), .B(n130), .C(n129), .D(\Queue[3][31] ), 
        .Z(n131) );
  OAI21M1P U308 ( .A(n206), .B(n132), .C(n131), .Z(n505) );
  OA21M1P U309 ( .A(n136), .B(n137), .C(Rst_n), .Z(n133) );
  AOI22M1P U310 ( .A(\Queue[3][0] ), .B(n203), .C(n202), .D(\Queue[4][0] ), 
        .Z(n140) );
  OAI21M1P U311 ( .A(n141), .B(n205), .C(n140), .Z(n506) );
  AOI22M1P U312 ( .A(\Queue[3][1] ), .B(n203), .C(n202), .D(\Queue[4][1] ), 
        .Z(n142) );
  OAI21M1P U313 ( .A(n143), .B(n205), .C(n142), .Z(n507) );
  AOI22M1P U314 ( .A(\Queue[3][2] ), .B(n203), .C(n202), .D(\Queue[4][2] ), 
        .Z(n144) );
  OAI21M1P U315 ( .A(n145), .B(n205), .C(n144), .Z(n508) );
  AOI22M1P U316 ( .A(\Queue[3][3] ), .B(n203), .C(n202), .D(\Queue[4][3] ), 
        .Z(n146) );
  OAI21M1P U317 ( .A(n147), .B(n205), .C(n146), .Z(n509) );
  AOI22M1P U318 ( .A(\Queue[3][4] ), .B(n203), .C(n202), .D(\Queue[4][4] ), 
        .Z(n148) );
  OAI21M1P U319 ( .A(n149), .B(n205), .C(n148), .Z(n510) );
  AOI22M1P U320 ( .A(\Queue[3][5] ), .B(n203), .C(n202), .D(\Queue[4][5] ), 
        .Z(n150) );
  OAI21M1P U321 ( .A(n151), .B(n205), .C(n150), .Z(n511) );
  AOI22M1P U322 ( .A(\Queue[3][6] ), .B(n203), .C(n202), .D(\Queue[4][6] ), 
        .Z(n152) );
  OAI21M1P U323 ( .A(n153), .B(n205), .C(n152), .Z(n512) );
  AOI22M1P U324 ( .A(\Queue[3][7] ), .B(n203), .C(n202), .D(\Queue[4][7] ), 
        .Z(n154) );
  OAI21M1P U325 ( .A(n155), .B(n205), .C(n154), .Z(n513) );
  AOI22M1P U326 ( .A(\Queue[3][8] ), .B(n203), .C(n202), .D(\Queue[4][8] ), 
        .Z(n156) );
  OAI21M1P U327 ( .A(n157), .B(n205), .C(n156), .Z(n514) );
  AOI22M1P U328 ( .A(\Queue[3][9] ), .B(n203), .C(n202), .D(\Queue[4][9] ), 
        .Z(n158) );
  OAI21M1P U329 ( .A(n159), .B(n205), .C(n158), .Z(n515) );
  AOI22M1P U330 ( .A(\Queue[3][10] ), .B(n203), .C(n202), .D(\Queue[4][10] ), 
        .Z(n160) );
  OAI21M1P U331 ( .A(n161), .B(n205), .C(n160), .Z(n516) );
  AOI22M1P U332 ( .A(\Queue[3][11] ), .B(n203), .C(n202), .D(\Queue[4][11] ), 
        .Z(n162) );
  OAI21M1P U333 ( .A(n163), .B(n205), .C(n162), .Z(n517) );
  AOI22M1P U334 ( .A(\Queue[3][12] ), .B(n203), .C(n202), .D(\Queue[4][12] ), 
        .Z(n164) );
  OAI21M1P U335 ( .A(n165), .B(n205), .C(n164), .Z(n518) );
  AOI22M1P U336 ( .A(\Queue[3][13] ), .B(n203), .C(n202), .D(\Queue[4][13] ), 
        .Z(n166) );
  OAI21M1P U337 ( .A(n167), .B(n205), .C(n166), .Z(n519) );
  AOI22M1P U338 ( .A(\Queue[3][14] ), .B(n203), .C(n202), .D(\Queue[4][14] ), 
        .Z(n168) );
  OAI21M1P U339 ( .A(n169), .B(n205), .C(n168), .Z(n520) );
  AOI22M1P U340 ( .A(\Queue[3][15] ), .B(n203), .C(n202), .D(\Queue[4][15] ), 
        .Z(n170) );
  OAI21M1P U341 ( .A(n171), .B(n205), .C(n170), .Z(n521) );
  AOI22M1P U342 ( .A(\Queue[3][16] ), .B(n203), .C(n202), .D(\Queue[4][16] ), 
        .Z(n172) );
  OAI21M1P U343 ( .A(n173), .B(n205), .C(n172), .Z(n522) );
  AOI22M1P U344 ( .A(\Queue[3][17] ), .B(n203), .C(n202), .D(\Queue[4][17] ), 
        .Z(n174) );
  OAI21M1P U345 ( .A(n175), .B(n205), .C(n174), .Z(n523) );
  AOI22M1P U346 ( .A(\Queue[3][18] ), .B(n203), .C(n202), .D(\Queue[4][18] ), 
        .Z(n176) );
  OAI21M1P U347 ( .A(n177), .B(n205), .C(n176), .Z(n524) );
  AOI22M1P U348 ( .A(\Queue[3][19] ), .B(n203), .C(n202), .D(\Queue[4][19] ), 
        .Z(n178) );
  OAI21M1P U349 ( .A(n179), .B(n205), .C(n178), .Z(n525) );
  AOI22M1P U350 ( .A(\Queue[3][20] ), .B(n203), .C(n202), .D(\Queue[4][20] ), 
        .Z(n180) );
  OAI21M1P U351 ( .A(n181), .B(n205), .C(n180), .Z(n526) );
  AOI22M1P U352 ( .A(\Queue[3][21] ), .B(n203), .C(n202), .D(\Queue[4][21] ), 
        .Z(n182) );
  OAI21M1P U353 ( .A(n183), .B(n205), .C(n182), .Z(n527) );
  AOI22M1P U354 ( .A(\Queue[3][22] ), .B(n203), .C(n202), .D(\Queue[4][22] ), 
        .Z(n184) );
  OAI21M1P U355 ( .A(n185), .B(n205), .C(n184), .Z(n528) );
  AOI22M1P U356 ( .A(\Queue[3][23] ), .B(n203), .C(n202), .D(\Queue[4][23] ), 
        .Z(n186) );
  OAI21M1P U357 ( .A(n187), .B(n205), .C(n186), .Z(n529) );
  AOI22M1P U358 ( .A(\Queue[3][24] ), .B(n203), .C(n202), .D(\Queue[4][24] ), 
        .Z(n188) );
  OAI21M1P U359 ( .A(n189), .B(n205), .C(n188), .Z(n530) );
  AOI22M1P U360 ( .A(\Queue[3][25] ), .B(n203), .C(n202), .D(\Queue[4][25] ), 
        .Z(n190) );
  OAI21M1P U361 ( .A(n191), .B(n205), .C(n190), .Z(n531) );
  AOI22M1P U362 ( .A(\Queue[3][26] ), .B(n203), .C(n202), .D(\Queue[4][26] ), 
        .Z(n192) );
  OAI21M1P U363 ( .A(n193), .B(n205), .C(n192), .Z(n532) );
  AOI22M1P U364 ( .A(\Queue[3][27] ), .B(n203), .C(n202), .D(\Queue[4][27] ), 
        .Z(n194) );
  OAI21M1P U365 ( .A(n195), .B(n205), .C(n194), .Z(n533) );
  AOI22M1P U366 ( .A(\Queue[3][28] ), .B(n203), .C(n202), .D(\Queue[4][28] ), 
        .Z(n196) );
  OAI21M1P U367 ( .A(n197), .B(n205), .C(n196), .Z(n534) );
  AOI22M1P U368 ( .A(\Queue[3][29] ), .B(n203), .C(n202), .D(\Queue[4][29] ), 
        .Z(n198) );
  OAI21M1P U369 ( .A(n199), .B(n205), .C(n198), .Z(n535) );
  AOI22M1P U370 ( .A(\Queue[3][30] ), .B(n203), .C(n202), .D(\Queue[4][30] ), 
        .Z(n200) );
  OAI21M1P U371 ( .A(n201), .B(n205), .C(n200), .Z(n536) );
  AOI22M1P U372 ( .A(\Queue[3][31] ), .B(n203), .C(n202), .D(\Queue[4][31] ), 
        .Z(n204) );
  OAI21M1P U373 ( .A(n206), .B(n205), .C(n204), .Z(n537) );
  N1M1P U374 ( .A(n538), .Z(Empty) );
  AOI22M1P U375 ( .A(n373), .B(n208), .C(n207), .D(Empty), .Z(n539) );
endmodule


module Packet_Queue_8 ( Clk_r, Rst_n, Packet_In, Read_Ack, Write_Ack, 
        Packet_Out, Empty, Full );
  input [31:0] Packet_In;
  output [31:0] Packet_Out;
  input Clk_r, Rst_n, Read_Ack, Write_Ack;
  output Empty, Full;
  wire   \Queue[4][31] , \Queue[4][30] , \Queue[4][29] , \Queue[4][28] ,
         \Queue[4][27] , \Queue[4][26] , \Queue[4][25] , \Queue[4][24] ,
         \Queue[4][23] , \Queue[4][22] , \Queue[4][21] , \Queue[4][20] ,
         \Queue[4][19] , \Queue[4][18] , \Queue[4][17] , \Queue[4][16] ,
         \Queue[4][15] , \Queue[4][14] , \Queue[4][13] , \Queue[4][12] ,
         \Queue[4][11] , \Queue[4][10] , \Queue[4][9] , \Queue[4][8] ,
         \Queue[4][7] , \Queue[4][6] , \Queue[4][5] , \Queue[4][4] ,
         \Queue[4][3] , \Queue[4][2] , \Queue[4][1] , \Queue[4][0] ,
         \Queue[3][31] , \Queue[3][30] , \Queue[3][29] , \Queue[3][28] ,
         \Queue[3][27] , \Queue[3][26] , \Queue[3][25] , \Queue[3][24] ,
         \Queue[3][23] , \Queue[3][22] , \Queue[3][21] , \Queue[3][20] ,
         \Queue[3][19] , \Queue[3][18] , \Queue[3][17] , \Queue[3][16] ,
         \Queue[3][15] , \Queue[3][14] , \Queue[3][13] , \Queue[3][12] ,
         \Queue[3][11] , \Queue[3][10] , \Queue[3][9] , \Queue[3][8] ,
         \Queue[3][7] , \Queue[3][6] , \Queue[3][5] , \Queue[3][4] ,
         \Queue[3][3] , \Queue[3][2] , \Queue[3][1] , \Queue[3][0] ,
         \Queue[2][31] , \Queue[2][30] , \Queue[2][29] , \Queue[2][28] ,
         \Queue[2][27] , \Queue[2][26] , \Queue[2][25] , \Queue[2][24] ,
         \Queue[2][23] , \Queue[2][22] , \Queue[2][21] , \Queue[2][20] ,
         \Queue[2][19] , \Queue[2][18] , \Queue[2][17] , \Queue[2][16] ,
         \Queue[2][15] , \Queue[2][14] , \Queue[2][13] , \Queue[2][12] ,
         \Queue[2][11] , \Queue[2][10] , \Queue[2][9] , \Queue[2][8] ,
         \Queue[2][7] , \Queue[2][6] , \Queue[2][5] , \Queue[2][4] ,
         \Queue[2][3] , \Queue[2][2] , \Queue[2][1] , \Queue[2][0] ,
         \Queue[1][31] , \Queue[1][30] , \Queue[1][29] , \Queue[1][28] ,
         \Queue[1][27] , \Queue[1][26] , \Queue[1][25] , \Queue[1][24] ,
         \Queue[1][23] , \Queue[1][22] , \Queue[1][21] , \Queue[1][20] ,
         \Queue[1][19] , \Queue[1][18] , \Queue[1][17] , \Queue[1][16] ,
         \Queue[1][15] , \Queue[1][14] , \Queue[1][13] , \Queue[1][12] ,
         \Queue[1][11] , \Queue[1][10] , \Queue[1][9] , \Queue[1][8] ,
         \Queue[1][7] , \Queue[1][6] , \Queue[1][5] , \Queue[1][4] ,
         \Queue[1][3] , \Queue[1][2] , \Queue[1][1] , \Queue[1][0] , n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541;
  wire   [2:0] Count;

  FDN2QM1P \Count_reg[0]  ( .D(n376), .CPN(Clk_r), .CD(Rst_n), .Q(Count[0]) );
  FDN2QM1P \Count_reg[1]  ( .D(n377), .CPN(Clk_r), .CD(Rst_n), .Q(Count[1]) );
  FDN2QM1P \Count_reg[2]  ( .D(n378), .CPN(Clk_r), .CD(Rst_n), .Q(Count[2]) );
  FDN1QM1P \Queue_reg[4][30]  ( .D(n410), .CPN(Clk_r), .Q(\Queue[4][30] ) );
  FDN1QM1P \Queue_reg[3][30]  ( .D(n538), .CPN(Clk_r), .Q(\Queue[3][30] ) );
  FDN1QM1P \Queue_reg[2][30]  ( .D(n506), .CPN(Clk_r), .Q(\Queue[2][30] ) );
  FDN1QM1P \Queue_reg[4][29]  ( .D(n409), .CPN(Clk_r), .Q(\Queue[4][29] ) );
  FDN1QM1P \Queue_reg[3][29]  ( .D(n537), .CPN(Clk_r), .Q(\Queue[3][29] ) );
  FDN1QM1P \Queue_reg[2][29]  ( .D(n505), .CPN(Clk_r), .Q(\Queue[2][29] ) );
  FDN1QM1P \Queue_reg[4][28]  ( .D(n408), .CPN(Clk_r), .Q(\Queue[4][28] ) );
  FDN1QM1P \Queue_reg[3][28]  ( .D(n536), .CPN(Clk_r), .Q(\Queue[3][28] ) );
  FDN1QM1P \Queue_reg[2][28]  ( .D(n504), .CPN(Clk_r), .Q(\Queue[2][28] ) );
  FDN1QM1P \Queue_reg[4][27]  ( .D(n407), .CPN(Clk_r), .Q(\Queue[4][27] ) );
  FDN1QM1P \Queue_reg[3][27]  ( .D(n535), .CPN(Clk_r), .Q(\Queue[3][27] ) );
  FDN1QM1P \Queue_reg[2][27]  ( .D(n503), .CPN(Clk_r), .Q(\Queue[2][27] ) );
  FDN1QM1P \Queue_reg[4][26]  ( .D(n406), .CPN(Clk_r), .Q(\Queue[4][26] ) );
  FDN1QM1P \Queue_reg[3][26]  ( .D(n534), .CPN(Clk_r), .Q(\Queue[3][26] ) );
  FDN1QM1P \Queue_reg[2][26]  ( .D(n502), .CPN(Clk_r), .Q(\Queue[2][26] ) );
  FDN1QM1P \Queue_reg[4][25]  ( .D(n405), .CPN(Clk_r), .Q(\Queue[4][25] ) );
  FDN1QM1P \Queue_reg[3][25]  ( .D(n533), .CPN(Clk_r), .Q(\Queue[3][25] ) );
  FDN1QM1P \Queue_reg[2][25]  ( .D(n501), .CPN(Clk_r), .Q(\Queue[2][25] ) );
  FDN1QM1P \Queue_reg[4][24]  ( .D(n404), .CPN(Clk_r), .Q(\Queue[4][24] ) );
  FDN1QM1P \Queue_reg[3][24]  ( .D(n532), .CPN(Clk_r), .Q(\Queue[3][24] ) );
  FDN1QM1P \Queue_reg[2][24]  ( .D(n500), .CPN(Clk_r), .Q(\Queue[2][24] ) );
  FDN1QM1P \Queue_reg[4][23]  ( .D(n403), .CPN(Clk_r), .Q(\Queue[4][23] ) );
  FDN1QM1P \Queue_reg[3][23]  ( .D(n531), .CPN(Clk_r), .Q(\Queue[3][23] ) );
  FDN1QM1P \Queue_reg[2][23]  ( .D(n499), .CPN(Clk_r), .Q(\Queue[2][23] ) );
  FDN1QM1P \Queue_reg[4][22]  ( .D(n402), .CPN(Clk_r), .Q(\Queue[4][22] ) );
  FDN1QM1P \Queue_reg[3][22]  ( .D(n530), .CPN(Clk_r), .Q(\Queue[3][22] ) );
  FDN1QM1P \Queue_reg[2][22]  ( .D(n498), .CPN(Clk_r), .Q(\Queue[2][22] ) );
  FDN1QM1P \Queue_reg[4][21]  ( .D(n401), .CPN(Clk_r), .Q(\Queue[4][21] ) );
  FDN1QM1P \Queue_reg[3][21]  ( .D(n529), .CPN(Clk_r), .Q(\Queue[3][21] ) );
  FDN1QM1P \Queue_reg[2][21]  ( .D(n497), .CPN(Clk_r), .Q(\Queue[2][21] ) );
  FDN1QM1P \Queue_reg[4][20]  ( .D(n400), .CPN(Clk_r), .Q(\Queue[4][20] ) );
  FDN1QM1P \Queue_reg[3][20]  ( .D(n528), .CPN(Clk_r), .Q(\Queue[3][20] ) );
  FDN1QM1P \Queue_reg[2][20]  ( .D(n496), .CPN(Clk_r), .Q(\Queue[2][20] ) );
  FDN1QM1P \Queue_reg[4][19]  ( .D(n399), .CPN(Clk_r), .Q(\Queue[4][19] ) );
  FDN1QM1P \Queue_reg[3][19]  ( .D(n527), .CPN(Clk_r), .Q(\Queue[3][19] ) );
  FDN1QM1P \Queue_reg[2][19]  ( .D(n495), .CPN(Clk_r), .Q(\Queue[2][19] ) );
  FDN1QM1P \Queue_reg[4][18]  ( .D(n398), .CPN(Clk_r), .Q(\Queue[4][18] ) );
  FDN1QM1P \Queue_reg[3][18]  ( .D(n526), .CPN(Clk_r), .Q(\Queue[3][18] ) );
  FDN1QM1P \Queue_reg[2][18]  ( .D(n494), .CPN(Clk_r), .Q(\Queue[2][18] ) );
  FDN1QM1P \Queue_reg[4][17]  ( .D(n397), .CPN(Clk_r), .Q(\Queue[4][17] ) );
  FDN1QM1P \Queue_reg[3][17]  ( .D(n525), .CPN(Clk_r), .Q(\Queue[3][17] ) );
  FDN1QM1P \Queue_reg[2][17]  ( .D(n493), .CPN(Clk_r), .Q(\Queue[2][17] ) );
  FDN1QM1P \Queue_reg[4][16]  ( .D(n396), .CPN(Clk_r), .Q(\Queue[4][16] ) );
  FDN1QM1P \Queue_reg[3][16]  ( .D(n524), .CPN(Clk_r), .Q(\Queue[3][16] ) );
  FDN1QM1P \Queue_reg[2][16]  ( .D(n492), .CPN(Clk_r), .Q(\Queue[2][16] ) );
  FDN1QM1P \Queue_reg[4][15]  ( .D(n395), .CPN(Clk_r), .Q(\Queue[4][15] ) );
  FDN1QM1P \Queue_reg[3][15]  ( .D(n523), .CPN(Clk_r), .Q(\Queue[3][15] ) );
  FDN1QM1P \Queue_reg[2][15]  ( .D(n491), .CPN(Clk_r), .Q(\Queue[2][15] ) );
  FDN1QM1P \Queue_reg[4][14]  ( .D(n394), .CPN(Clk_r), .Q(\Queue[4][14] ) );
  FDN1QM1P \Queue_reg[3][14]  ( .D(n522), .CPN(Clk_r), .Q(\Queue[3][14] ) );
  FDN1QM1P \Queue_reg[2][14]  ( .D(n490), .CPN(Clk_r), .Q(\Queue[2][14] ) );
  FDN1QM1P \Queue_reg[4][13]  ( .D(n393), .CPN(Clk_r), .Q(\Queue[4][13] ) );
  FDN1QM1P \Queue_reg[3][13]  ( .D(n521), .CPN(Clk_r), .Q(\Queue[3][13] ) );
  FDN1QM1P \Queue_reg[2][13]  ( .D(n489), .CPN(Clk_r), .Q(\Queue[2][13] ) );
  FDN1QM1P \Queue_reg[4][12]  ( .D(n392), .CPN(Clk_r), .Q(\Queue[4][12] ) );
  FDN1QM1P \Queue_reg[3][12]  ( .D(n520), .CPN(Clk_r), .Q(\Queue[3][12] ) );
  FDN1QM1P \Queue_reg[2][12]  ( .D(n488), .CPN(Clk_r), .Q(\Queue[2][12] ) );
  FDN1QM1P \Queue_reg[4][11]  ( .D(n391), .CPN(Clk_r), .Q(\Queue[4][11] ) );
  FDN1QM1P \Queue_reg[3][11]  ( .D(n519), .CPN(Clk_r), .Q(\Queue[3][11] ) );
  FDN1QM1P \Queue_reg[2][11]  ( .D(n487), .CPN(Clk_r), .Q(\Queue[2][11] ) );
  FDN1QM1P \Queue_reg[4][10]  ( .D(n390), .CPN(Clk_r), .Q(\Queue[4][10] ) );
  FDN1QM1P \Queue_reg[3][10]  ( .D(n518), .CPN(Clk_r), .Q(\Queue[3][10] ) );
  FDN1QM1P \Queue_reg[2][10]  ( .D(n486), .CPN(Clk_r), .Q(\Queue[2][10] ) );
  FDN1QM1P \Queue_reg[4][9]  ( .D(n389), .CPN(Clk_r), .Q(\Queue[4][9] ) );
  FDN1QM1P \Queue_reg[3][9]  ( .D(n517), .CPN(Clk_r), .Q(\Queue[3][9] ) );
  FDN1QM1P \Queue_reg[2][9]  ( .D(n485), .CPN(Clk_r), .Q(\Queue[2][9] ) );
  FDN1QM1P \Queue_reg[4][8]  ( .D(n388), .CPN(Clk_r), .Q(\Queue[4][8] ) );
  FDN1QM1P \Queue_reg[3][8]  ( .D(n516), .CPN(Clk_r), .Q(\Queue[3][8] ) );
  FDN1QM1P \Queue_reg[2][8]  ( .D(n484), .CPN(Clk_r), .Q(\Queue[2][8] ) );
  FDN1QM1P \Queue_reg[4][7]  ( .D(n387), .CPN(Clk_r), .Q(\Queue[4][7] ) );
  FDN1QM1P \Queue_reg[3][7]  ( .D(n515), .CPN(Clk_r), .Q(\Queue[3][7] ) );
  FDN1QM1P \Queue_reg[2][7]  ( .D(n483), .CPN(Clk_r), .Q(\Queue[2][7] ) );
  FDN1QM1P \Queue_reg[4][6]  ( .D(n386), .CPN(Clk_r), .Q(\Queue[4][6] ) );
  FDN1QM1P \Queue_reg[3][6]  ( .D(n514), .CPN(Clk_r), .Q(\Queue[3][6] ) );
  FDN1QM1P \Queue_reg[2][6]  ( .D(n482), .CPN(Clk_r), .Q(\Queue[2][6] ) );
  FDN1QM1P \Queue_reg[4][5]  ( .D(n385), .CPN(Clk_r), .Q(\Queue[4][5] ) );
  FDN1QM1P \Queue_reg[3][5]  ( .D(n513), .CPN(Clk_r), .Q(\Queue[3][5] ) );
  FDN1QM1P \Queue_reg[2][5]  ( .D(n481), .CPN(Clk_r), .Q(\Queue[2][5] ) );
  FDN1QM1P \Queue_reg[4][4]  ( .D(n384), .CPN(Clk_r), .Q(\Queue[4][4] ) );
  FDN1QM1P \Queue_reg[3][4]  ( .D(n512), .CPN(Clk_r), .Q(\Queue[3][4] ) );
  FDN1QM1P \Queue_reg[2][4]  ( .D(n480), .CPN(Clk_r), .Q(\Queue[2][4] ) );
  FDN1QM1P \Queue_reg[4][3]  ( .D(n383), .CPN(Clk_r), .Q(\Queue[4][3] ) );
  FDN1QM1P \Queue_reg[3][3]  ( .D(n511), .CPN(Clk_r), .Q(\Queue[3][3] ) );
  FDN1QM1P \Queue_reg[2][3]  ( .D(n479), .CPN(Clk_r), .Q(\Queue[2][3] ) );
  FDN1QM1P \Queue_reg[4][2]  ( .D(n382), .CPN(Clk_r), .Q(\Queue[4][2] ) );
  FDN1QM1P \Queue_reg[3][2]  ( .D(n510), .CPN(Clk_r), .Q(\Queue[3][2] ) );
  FDN1QM1P \Queue_reg[2][2]  ( .D(n478), .CPN(Clk_r), .Q(\Queue[2][2] ) );
  FDN1QM1P \Queue_reg[4][1]  ( .D(n381), .CPN(Clk_r), .Q(\Queue[4][1] ) );
  FDN1QM1P \Queue_reg[3][1]  ( .D(n509), .CPN(Clk_r), .Q(\Queue[3][1] ) );
  FDN1QM1P \Queue_reg[2][1]  ( .D(n477), .CPN(Clk_r), .Q(\Queue[2][1] ) );
  FDN1QM1P \Queue_reg[4][0]  ( .D(n380), .CPN(Clk_r), .Q(\Queue[4][0] ) );
  FDN1QM1P \Queue_reg[3][0]  ( .D(n508), .CPN(Clk_r), .Q(\Queue[3][0] ) );
  FDN1QM1P \Queue_reg[2][0]  ( .D(n476), .CPN(Clk_r), .Q(\Queue[2][0] ) );
  FDN1QM1P \Queue_reg[4][31]  ( .D(n379), .CPN(Clk_r), .Q(\Queue[4][31] ) );
  FDN1QM1P \Queue_reg[3][31]  ( .D(n539), .CPN(Clk_r), .Q(\Queue[3][31] ) );
  FDN1QM1P \Queue_reg[2][31]  ( .D(n507), .CPN(Clk_r), .Q(\Queue[2][31] ) );
  FDN2QM1P Full_reg ( .D(n411), .CPN(Clk_r), .CD(Rst_n), .Q(Full) );
  FDN1QM1P \Queue_reg[1][31]  ( .D(n443), .CPN(Clk_r), .Q(\Queue[1][31] ) );
  FDN1QM1P \Queue_reg[0][31]  ( .D(n475), .CPN(Clk_r), .Q(Packet_Out[31]) );
  FDN1QM1P \Queue_reg[1][30]  ( .D(n442), .CPN(Clk_r), .Q(\Queue[1][30] ) );
  FDN1QM1P \Queue_reg[0][30]  ( .D(n474), .CPN(Clk_r), .Q(Packet_Out[30]) );
  FDN1QM1P \Queue_reg[1][29]  ( .D(n441), .CPN(Clk_r), .Q(\Queue[1][29] ) );
  FDN1QM1P \Queue_reg[0][29]  ( .D(n473), .CPN(Clk_r), .Q(Packet_Out[29]) );
  FDN1QM1P \Queue_reg[1][28]  ( .D(n440), .CPN(Clk_r), .Q(\Queue[1][28] ) );
  FDN1QM1P \Queue_reg[0][28]  ( .D(n472), .CPN(Clk_r), .Q(Packet_Out[28]) );
  FDN1QM1P \Queue_reg[1][27]  ( .D(n439), .CPN(Clk_r), .Q(\Queue[1][27] ) );
  FDN1QM1P \Queue_reg[0][27]  ( .D(n471), .CPN(Clk_r), .Q(Packet_Out[27]) );
  FDN1QM1P \Queue_reg[1][26]  ( .D(n438), .CPN(Clk_r), .Q(\Queue[1][26] ) );
  FDN1QM1P \Queue_reg[0][26]  ( .D(n470), .CPN(Clk_r), .Q(Packet_Out[26]) );
  FDN1QM1P \Queue_reg[1][25]  ( .D(n437), .CPN(Clk_r), .Q(\Queue[1][25] ) );
  FDN1QM1P \Queue_reg[0][25]  ( .D(n469), .CPN(Clk_r), .Q(Packet_Out[25]) );
  FDN1QM1P \Queue_reg[1][24]  ( .D(n436), .CPN(Clk_r), .Q(\Queue[1][24] ) );
  FDN1QM1P \Queue_reg[0][24]  ( .D(n468), .CPN(Clk_r), .Q(Packet_Out[24]) );
  FDN1QM1P \Queue_reg[1][23]  ( .D(n435), .CPN(Clk_r), .Q(\Queue[1][23] ) );
  FDN1QM1P \Queue_reg[0][23]  ( .D(n467), .CPN(Clk_r), .Q(Packet_Out[23]) );
  FDN1QM1P \Queue_reg[1][22]  ( .D(n434), .CPN(Clk_r), .Q(\Queue[1][22] ) );
  FDN1QM1P \Queue_reg[0][22]  ( .D(n466), .CPN(Clk_r), .Q(Packet_Out[22]) );
  FDN1QM1P \Queue_reg[1][21]  ( .D(n433), .CPN(Clk_r), .Q(\Queue[1][21] ) );
  FDN1QM1P \Queue_reg[0][21]  ( .D(n465), .CPN(Clk_r), .Q(Packet_Out[21]) );
  FDN1QM1P \Queue_reg[1][20]  ( .D(n432), .CPN(Clk_r), .Q(\Queue[1][20] ) );
  FDN1QM1P \Queue_reg[0][20]  ( .D(n464), .CPN(Clk_r), .Q(Packet_Out[20]) );
  FDN1QM1P \Queue_reg[1][19]  ( .D(n431), .CPN(Clk_r), .Q(\Queue[1][19] ) );
  FDN1QM1P \Queue_reg[0][19]  ( .D(n463), .CPN(Clk_r), .Q(Packet_Out[19]) );
  FDN1QM1P \Queue_reg[1][18]  ( .D(n430), .CPN(Clk_r), .Q(\Queue[1][18] ) );
  FDN1QM1P \Queue_reg[0][18]  ( .D(n462), .CPN(Clk_r), .Q(Packet_Out[18]) );
  FDN1QM1P \Queue_reg[1][17]  ( .D(n429), .CPN(Clk_r), .Q(\Queue[1][17] ) );
  FDN1QM1P \Queue_reg[0][17]  ( .D(n461), .CPN(Clk_r), .Q(Packet_Out[17]) );
  FDN1QM1P \Queue_reg[1][16]  ( .D(n428), .CPN(Clk_r), .Q(\Queue[1][16] ) );
  FDN1QM1P \Queue_reg[0][16]  ( .D(n460), .CPN(Clk_r), .Q(Packet_Out[16]) );
  FDN1QM1P \Queue_reg[1][15]  ( .D(n427), .CPN(Clk_r), .Q(\Queue[1][15] ) );
  FDN1QM1P \Queue_reg[0][15]  ( .D(n459), .CPN(Clk_r), .Q(Packet_Out[15]) );
  FDN1QM1P \Queue_reg[1][14]  ( .D(n426), .CPN(Clk_r), .Q(\Queue[1][14] ) );
  FDN1QM1P \Queue_reg[0][14]  ( .D(n458), .CPN(Clk_r), .Q(Packet_Out[14]) );
  FDN1QM1P \Queue_reg[1][13]  ( .D(n425), .CPN(Clk_r), .Q(\Queue[1][13] ) );
  FDN1QM1P \Queue_reg[0][13]  ( .D(n457), .CPN(Clk_r), .Q(Packet_Out[13]) );
  FDN1QM1P \Queue_reg[1][12]  ( .D(n424), .CPN(Clk_r), .Q(\Queue[1][12] ) );
  FDN1QM1P \Queue_reg[0][12]  ( .D(n456), .CPN(Clk_r), .Q(Packet_Out[12]) );
  FDN1QM1P \Queue_reg[1][11]  ( .D(n423), .CPN(Clk_r), .Q(\Queue[1][11] ) );
  FDN1QM1P \Queue_reg[0][11]  ( .D(n455), .CPN(Clk_r), .Q(Packet_Out[11]) );
  FDN1QM1P \Queue_reg[1][10]  ( .D(n422), .CPN(Clk_r), .Q(\Queue[1][10] ) );
  FDN1QM1P \Queue_reg[0][10]  ( .D(n454), .CPN(Clk_r), .Q(Packet_Out[10]) );
  FDN1QM1P \Queue_reg[1][9]  ( .D(n421), .CPN(Clk_r), .Q(\Queue[1][9] ) );
  FDN1QM1P \Queue_reg[0][9]  ( .D(n453), .CPN(Clk_r), .Q(Packet_Out[9]) );
  FDN1QM1P \Queue_reg[1][8]  ( .D(n420), .CPN(Clk_r), .Q(\Queue[1][8] ) );
  FDN1QM1P \Queue_reg[0][8]  ( .D(n452), .CPN(Clk_r), .Q(Packet_Out[8]) );
  FDN1QM1P \Queue_reg[1][7]  ( .D(n419), .CPN(Clk_r), .Q(\Queue[1][7] ) );
  FDN1QM1P \Queue_reg[0][7]  ( .D(n451), .CPN(Clk_r), .Q(Packet_Out[7]) );
  FDN1QM1P \Queue_reg[1][6]  ( .D(n418), .CPN(Clk_r), .Q(\Queue[1][6] ) );
  FDN1QM1P \Queue_reg[0][6]  ( .D(n450), .CPN(Clk_r), .Q(Packet_Out[6]) );
  FDN1QM1P \Queue_reg[1][5]  ( .D(n417), .CPN(Clk_r), .Q(\Queue[1][5] ) );
  FDN1QM1P \Queue_reg[0][5]  ( .D(n449), .CPN(Clk_r), .Q(Packet_Out[5]) );
  FDN1QM1P \Queue_reg[1][4]  ( .D(n416), .CPN(Clk_r), .Q(\Queue[1][4] ) );
  FDN1QM1P \Queue_reg[0][4]  ( .D(n448), .CPN(Clk_r), .Q(Packet_Out[4]) );
  FDN1QM1P \Queue_reg[1][3]  ( .D(n415), .CPN(Clk_r), .Q(\Queue[1][3] ) );
  FDN1QM1P \Queue_reg[0][3]  ( .D(n447), .CPN(Clk_r), .Q(Packet_Out[3]) );
  FDN1QM1P \Queue_reg[1][2]  ( .D(n414), .CPN(Clk_r), .Q(\Queue[1][2] ) );
  FDN1QM1P \Queue_reg[0][2]  ( .D(n446), .CPN(Clk_r), .Q(Packet_Out[2]) );
  FDN1QM1P \Queue_reg[1][1]  ( .D(n413), .CPN(Clk_r), .Q(\Queue[1][1] ) );
  FDN1QM1P \Queue_reg[0][1]  ( .D(n445), .CPN(Clk_r), .Q(Packet_Out[1]) );
  FDN1QM1P \Queue_reg[1][0]  ( .D(n412), .CPN(Clk_r), .Q(\Queue[1][0] ) );
  FDN1QM1P \Queue_reg[0][0]  ( .D(n444), .CPN(Clk_r), .Q(Packet_Out[0]) );
  FDN2QM1P Empty_reg ( .D(n541), .CPN(Clk_r), .CD(Rst_n), .Q(n540) );
  BUFM2P U3 ( .A(n58), .Z(n7) );
  BUFM2P U4 ( .A(n96), .Z(n8) );
  BUFM1P U5 ( .A(n96), .Z(n9) );
  BUFM1P U6 ( .A(n205), .Z(n11) );
  BUFM2P U7 ( .A(n205), .Z(n10) );
  N1M1P U8 ( .A(Read_Ack), .Z(n136) );
  BUFM3P U9 ( .A(n55), .Z(n5) );
  AOI21M3P U10 ( .A(n3), .B(n99), .C(n140), .Z(n56) );
  AOI21M3P U11 ( .A(n3), .B(n141), .C(n140), .Z(n204) );
  AOI21M3P U12 ( .A(n3), .B(n139), .C(n140), .Z(n131) );
  OAI211M4P U13 ( .A(n139), .B(n136), .C(n3), .D(n97), .Z(n134) );
  OAI211M4P U14 ( .A(n141), .B(n136), .C(n3), .D(n135), .Z(n207) );
  NR2I1M8P U15 ( .A(n60), .B(n20), .Z(n19) );
  OAI211M4P U16 ( .A(n99), .B(n138), .C(Rst_n), .D(n137), .Z(n132) );
  N1M2P U17 ( .A(n61), .Z(n93) );
  OAI21M2P U18 ( .A(n3), .B(Read_Ack), .C(n23), .Z(n55) );
  BUFM2P U19 ( .A(n58), .Z(n6) );
  NR3M1P U20 ( .A(Count[2]), .B(n22), .C(n21), .Z(n139) );
  OAI211M2P U21 ( .A(n99), .B(n136), .C(n3), .D(n23), .Z(n58) );
  ND2M1P U22 ( .A(n17), .B(Rst_n), .Z(n60) );
  NR2FM1P U23 ( .A(Read_Ack), .B(n98), .Z(n17) );
  NR3M1P U24 ( .A(Count[0]), .B(Count[2]), .C(n21), .Z(n99) );
  NR3M1P U25 ( .A(Count[0]), .B(Count[1]), .C(n18), .Z(n141) );
  NR3M1P U26 ( .A(n22), .B(Count[2]), .C(Count[1]), .Z(n375) );
  N1M3P U27 ( .A(n3), .Z(n98) );
  N1M1P U28 ( .A(Count[1]), .Z(n21) );
  BUFM8P U29 ( .A(Write_Ack), .Z(n3) );
  N1M1P U30 ( .A(Count[0]), .Z(n22) );
  N1M1P U31 ( .A(Count[2]), .Z(n18) );
  N1M1P U32 ( .A(Packet_In[29]), .Z(n201) );
  N1M1P U33 ( .A(Packet_In[28]), .Z(n199) );
  N1M1P U34 ( .A(Packet_In[26]), .Z(n195) );
  N1M1P U35 ( .A(Packet_In[27]), .Z(n197) );
  N1M1P U36 ( .A(Packet_In[31]), .Z(n208) );
  N1M1P U37 ( .A(Packet_In[22]), .Z(n187) );
  N1M1P U38 ( .A(Packet_In[24]), .Z(n191) );
  N1M1P U39 ( .A(Packet_In[25]), .Z(n193) );
  N1M1P U40 ( .A(Packet_In[20]), .Z(n183) );
  N1M1P U41 ( .A(Packet_In[21]), .Z(n185) );
  N1M1P U42 ( .A(Packet_In[23]), .Z(n189) );
  N1M1P U43 ( .A(Packet_In[30]), .Z(n203) );
  N1M1P U44 ( .A(Packet_In[3]), .Z(n149) );
  N1M1P U45 ( .A(Packet_In[1]), .Z(n145) );
  N1M1P U46 ( .A(Packet_In[6]), .Z(n155) );
  N1M1P U47 ( .A(Packet_In[7]), .Z(n157) );
  N1M1P U48 ( .A(Packet_In[5]), .Z(n153) );
  N1M1P U49 ( .A(Packet_In[4]), .Z(n151) );
  N1M1P U50 ( .A(Packet_In[8]), .Z(n159) );
  N1M1P U51 ( .A(Packet_In[0]), .Z(n143) );
  N1M1P U52 ( .A(Packet_In[9]), .Z(n161) );
  N1M1P U53 ( .A(Packet_In[19]), .Z(n181) );
  N1M1P U54 ( .A(Packet_In[18]), .Z(n179) );
  N1M1P U55 ( .A(Packet_In[10]), .Z(n163) );
  N1M1P U56 ( .A(Packet_In[17]), .Z(n177) );
  N1M1P U57 ( .A(Packet_In[2]), .Z(n147) );
  N1M1P U58 ( .A(Packet_In[16]), .Z(n175) );
  N1M1P U59 ( .A(Packet_In[15]), .Z(n173) );
  N1M1P U60 ( .A(Packet_In[11]), .Z(n165) );
  N1M1P U61 ( .A(Packet_In[14]), .Z(n171) );
  N1M1P U62 ( .A(Packet_In[13]), .Z(n169) );
  N1M1P U63 ( .A(Packet_In[12]), .Z(n167) );
  BUFM2P U64 ( .A(n55), .Z(n4) );
  N1M2P U65 ( .A(n17), .Z(n138) );
  AOI21M6P U66 ( .A(n3), .B(n375), .C(n140), .Z(n94) );
  OAI211M1P U67 ( .A(n375), .B(n136), .C(n3), .D(n61), .Z(n96) );
  ND2M1P U68 ( .A(Read_Ack), .B(Rst_n), .Z(n140) );
  OAI211M1P U69 ( .A(n139), .B(n138), .C(Rst_n), .D(n137), .Z(n205) );
  NR2M1P U70 ( .A(n136), .B(n3), .Z(n374) );
  NR2M1P U71 ( .A(n17), .B(n374), .Z(n373) );
  AOI22CDNM1P U72 ( .A(n373), .B(n22), .C(n373), .D(n22), .Z(n376) );
  N1M1P U73 ( .A(n374), .Z(n16) );
  AOI22M1P U74 ( .A(Count[0]), .B(n138), .C(n16), .D(n22), .Z(n13) );
  AOI22CDNM1P U75 ( .A(Count[1]), .B(n13), .C(n13), .D(Count[1]), .Z(n377) );
  ND3M1P U76 ( .A(n22), .B(n18), .C(n21), .Z(n59) );
  ND2M1P U77 ( .A(Count[1]), .B(Read_Ack), .Z(n12) );
  OAI211M1P U78 ( .A(Count[1]), .B(n138), .C(n13), .D(n12), .Z(n14) );
  AOI22M1P U79 ( .A(n17), .B(n139), .C(Count[2]), .D(n14), .Z(n15) );
  OAI21M1P U80 ( .A(n59), .B(n16), .C(n15), .Z(n378) );
  N1M1P U81 ( .A(n141), .Z(n20) );
  AOI22CDNM1P U82 ( .A(n19), .B(n208), .C(\Queue[4][31] ), .D(n19), .Z(n379)
         );
  AOI22CDNM1P U83 ( .A(n19), .B(n143), .C(\Queue[4][0] ), .D(n19), .Z(n380) );
  AOI22CDNM1P U84 ( .A(n19), .B(n145), .C(\Queue[4][1] ), .D(n19), .Z(n381) );
  AOI22CDNM1P U85 ( .A(n19), .B(n147), .C(\Queue[4][2] ), .D(n19), .Z(n382) );
  AOI22CDNM1P U86 ( .A(n19), .B(n149), .C(\Queue[4][3] ), .D(n19), .Z(n383) );
  AOI22CDNM1P U87 ( .A(n19), .B(n151), .C(\Queue[4][4] ), .D(n19), .Z(n384) );
  AOI22CDNM1P U88 ( .A(n19), .B(n153), .C(\Queue[4][5] ), .D(n19), .Z(n385) );
  AOI22CDNM1P U89 ( .A(n19), .B(n155), .C(\Queue[4][6] ), .D(n19), .Z(n386) );
  AOI22CDNM1P U90 ( .A(n19), .B(n157), .C(\Queue[4][7] ), .D(n19), .Z(n387) );
  AOI22CDNM1P U91 ( .A(n19), .B(n159), .C(\Queue[4][8] ), .D(n19), .Z(n388) );
  AOI22CDNM1P U92 ( .A(n19), .B(n161), .C(\Queue[4][9] ), .D(n19), .Z(n389) );
  AOI22CDNM1P U93 ( .A(n19), .B(n163), .C(\Queue[4][10] ), .D(n19), .Z(n390)
         );
  AOI22CDNM1P U94 ( .A(n19), .B(n165), .C(\Queue[4][11] ), .D(n19), .Z(n391)
         );
  AOI22CDNM1P U95 ( .A(n19), .B(n167), .C(\Queue[4][12] ), .D(n19), .Z(n392)
         );
  AOI22CDNM1P U96 ( .A(n19), .B(n169), .C(\Queue[4][13] ), .D(n19), .Z(n393)
         );
  AOI22CDNM1P U97 ( .A(n19), .B(n171), .C(\Queue[4][14] ), .D(n19), .Z(n394)
         );
  AOI22CDNM1P U98 ( .A(n19), .B(n173), .C(\Queue[4][15] ), .D(n19), .Z(n395)
         );
  AOI22CDNM1P U99 ( .A(n19), .B(n175), .C(\Queue[4][16] ), .D(n19), .Z(n396)
         );
  AOI22CDNM1P U100 ( .A(n19), .B(n177), .C(\Queue[4][17] ), .D(n19), .Z(n397)
         );
  AOI22CDNM1P U101 ( .A(n19), .B(n179), .C(\Queue[4][18] ), .D(n19), .Z(n398)
         );
  AOI22CDNM1P U102 ( .A(n19), .B(n181), .C(\Queue[4][19] ), .D(n19), .Z(n399)
         );
  AOI22CDNM1P U103 ( .A(n19), .B(n183), .C(\Queue[4][20] ), .D(n19), .Z(n400)
         );
  AOI22CDNM1P U104 ( .A(n19), .B(n185), .C(\Queue[4][21] ), .D(n19), .Z(n401)
         );
  AOI22CDNM1P U105 ( .A(n19), .B(n187), .C(\Queue[4][22] ), .D(n19), .Z(n402)
         );
  AOI22CDNM1P U106 ( .A(n19), .B(n189), .C(\Queue[4][23] ), .D(n19), .Z(n403)
         );
  AOI22CDNM1P U107 ( .A(n19), .B(n191), .C(\Queue[4][24] ), .D(n19), .Z(n404)
         );
  AOI22CDNM1P U108 ( .A(n19), .B(n193), .C(\Queue[4][25] ), .D(n19), .Z(n405)
         );
  AOI22CDNM1P U109 ( .A(n19), .B(n195), .C(\Queue[4][26] ), .D(n19), .Z(n406)
         );
  AOI22CDNM1P U110 ( .A(n19), .B(n197), .C(\Queue[4][27] ), .D(n19), .Z(n407)
         );
  AOI22CDNM1P U111 ( .A(n19), .B(n199), .C(\Queue[4][28] ), .D(n19), .Z(n408)
         );
  AOI22CDNM1P U112 ( .A(n19), .B(n201), .C(\Queue[4][29] ), .D(n19), .Z(n409)
         );
  AOI22CDNM1P U113 ( .A(n19), .B(n203), .C(\Queue[4][30] ), .D(n19), .Z(n410)
         );
  OAI22CDNM1P U114 ( .A(n138), .B(n20), .C(n373), .D(Full), .Z(n411) );
  OA21M1P U115 ( .A(n138), .B(n375), .C(Rst_n), .Z(n23) );
  AOI22M1P U116 ( .A(\Queue[2][0] ), .B(n56), .C(\Queue[1][0] ), .D(n4), .Z(
        n24) );
  OAI21M1P U117 ( .A(n143), .B(n7), .C(n24), .Z(n412) );
  AOI22M1P U118 ( .A(n56), .B(\Queue[2][1] ), .C(\Queue[1][1] ), .D(n4), .Z(
        n25) );
  OAI21M1P U119 ( .A(n6), .B(n145), .C(n25), .Z(n413) );
  AOI22M1P U120 ( .A(n56), .B(\Queue[2][2] ), .C(\Queue[1][2] ), .D(n4), .Z(
        n26) );
  OAI21M1P U121 ( .A(n7), .B(n147), .C(n26), .Z(n414) );
  AOI22M1P U122 ( .A(n56), .B(\Queue[2][3] ), .C(\Queue[1][3] ), .D(n4), .Z(
        n27) );
  OAI21M1P U123 ( .A(n7), .B(n149), .C(n27), .Z(n415) );
  AOI22M1P U124 ( .A(n56), .B(\Queue[2][4] ), .C(\Queue[1][4] ), .D(n4), .Z(
        n28) );
  OAI21M1P U125 ( .A(n7), .B(n151), .C(n28), .Z(n416) );
  AOI22M1P U126 ( .A(n56), .B(\Queue[2][5] ), .C(\Queue[1][5] ), .D(n4), .Z(
        n29) );
  OAI21M1P U127 ( .A(n7), .B(n153), .C(n29), .Z(n417) );
  AOI22M1P U128 ( .A(n56), .B(\Queue[2][6] ), .C(\Queue[1][6] ), .D(n4), .Z(
        n30) );
  OAI21M1P U129 ( .A(n7), .B(n155), .C(n30), .Z(n418) );
  AOI22M1P U130 ( .A(n56), .B(\Queue[2][7] ), .C(\Queue[1][7] ), .D(n4), .Z(
        n31) );
  OAI21M1P U131 ( .A(n7), .B(n157), .C(n31), .Z(n419) );
  AOI22M1P U132 ( .A(n56), .B(\Queue[2][8] ), .C(\Queue[1][8] ), .D(n4), .Z(
        n32) );
  OAI21M1P U133 ( .A(n7), .B(n159), .C(n32), .Z(n420) );
  AOI22M1P U134 ( .A(n56), .B(\Queue[2][9] ), .C(\Queue[1][9] ), .D(n55), .Z(
        n33) );
  OAI21M1P U135 ( .A(n7), .B(n161), .C(n33), .Z(n421) );
  AOI22M1P U136 ( .A(n56), .B(\Queue[2][10] ), .C(\Queue[1][10] ), .D(n55), 
        .Z(n34) );
  OAI21M1P U137 ( .A(n7), .B(n163), .C(n34), .Z(n422) );
  AOI22M1P U138 ( .A(n56), .B(\Queue[2][11] ), .C(\Queue[1][11] ), .D(n55), 
        .Z(n35) );
  OAI21M1P U139 ( .A(n7), .B(n165), .C(n35), .Z(n423) );
  AOI22M1P U140 ( .A(n56), .B(\Queue[2][12] ), .C(\Queue[1][12] ), .D(n55), 
        .Z(n36) );
  OAI21M1P U141 ( .A(n6), .B(n167), .C(n36), .Z(n424) );
  AOI22M1P U142 ( .A(n56), .B(\Queue[2][13] ), .C(\Queue[1][13] ), .D(n55), 
        .Z(n37) );
  OAI21M1P U143 ( .A(n6), .B(n169), .C(n37), .Z(n425) );
  AOI22M1P U144 ( .A(n56), .B(\Queue[2][14] ), .C(\Queue[1][14] ), .D(n55), 
        .Z(n38) );
  OAI21M1P U145 ( .A(n6), .B(n171), .C(n38), .Z(n426) );
  AOI22M1P U146 ( .A(n56), .B(\Queue[2][15] ), .C(\Queue[1][15] ), .D(n55), 
        .Z(n39) );
  OAI21M1P U147 ( .A(n6), .B(n173), .C(n39), .Z(n427) );
  AOI22M1P U148 ( .A(n56), .B(\Queue[2][16] ), .C(\Queue[1][16] ), .D(n5), .Z(
        n40) );
  OAI21M1P U149 ( .A(n6), .B(n175), .C(n40), .Z(n428) );
  AOI22M1P U150 ( .A(n56), .B(\Queue[2][17] ), .C(\Queue[1][17] ), .D(n4), .Z(
        n41) );
  OAI21M1P U151 ( .A(n6), .B(n177), .C(n41), .Z(n429) );
  AOI22M1P U152 ( .A(n56), .B(\Queue[2][18] ), .C(\Queue[1][18] ), .D(n5), .Z(
        n42) );
  OAI21M1P U153 ( .A(n6), .B(n179), .C(n42), .Z(n430) );
  AOI22M1P U154 ( .A(n56), .B(\Queue[2][19] ), .C(\Queue[1][19] ), .D(n5), .Z(
        n43) );
  OAI21M1P U155 ( .A(n6), .B(n181), .C(n43), .Z(n431) );
  AOI22M1P U156 ( .A(n56), .B(\Queue[2][20] ), .C(\Queue[1][20] ), .D(n5), .Z(
        n44) );
  OAI21M1P U157 ( .A(n6), .B(n183), .C(n44), .Z(n432) );
  AOI22M1P U158 ( .A(n56), .B(\Queue[2][21] ), .C(\Queue[1][21] ), .D(n5), .Z(
        n45) );
  OAI21M1P U159 ( .A(n6), .B(n185), .C(n45), .Z(n433) );
  AOI22M1P U160 ( .A(n56), .B(\Queue[2][22] ), .C(\Queue[1][22] ), .D(n5), .Z(
        n46) );
  OAI21M1P U161 ( .A(n7), .B(n187), .C(n46), .Z(n434) );
  AOI22M1P U162 ( .A(n56), .B(\Queue[2][23] ), .C(\Queue[1][23] ), .D(n5), .Z(
        n47) );
  OAI21M1P U163 ( .A(n6), .B(n189), .C(n47), .Z(n435) );
  AOI22M1P U164 ( .A(n56), .B(\Queue[2][24] ), .C(\Queue[1][24] ), .D(n5), .Z(
        n48) );
  OAI21M1P U165 ( .A(n7), .B(n191), .C(n48), .Z(n436) );
  AOI22M1P U166 ( .A(n56), .B(\Queue[2][25] ), .C(\Queue[1][25] ), .D(n5), .Z(
        n49) );
  OAI21M1P U167 ( .A(n6), .B(n193), .C(n49), .Z(n437) );
  AOI22M1P U168 ( .A(n56), .B(\Queue[2][26] ), .C(\Queue[1][26] ), .D(n5), .Z(
        n50) );
  OAI21M1P U169 ( .A(n58), .B(n195), .C(n50), .Z(n438) );
  AOI22M1P U170 ( .A(n56), .B(\Queue[2][27] ), .C(\Queue[1][27] ), .D(n5), .Z(
        n51) );
  OAI21M1P U171 ( .A(n58), .B(n197), .C(n51), .Z(n439) );
  AOI22M1P U172 ( .A(n56), .B(\Queue[2][28] ), .C(\Queue[1][28] ), .D(n4), .Z(
        n52) );
  OAI21M1P U173 ( .A(n58), .B(n199), .C(n52), .Z(n440) );
  AOI22M1P U174 ( .A(n56), .B(\Queue[2][29] ), .C(\Queue[1][29] ), .D(n5), .Z(
        n53) );
  OAI21M1P U175 ( .A(n58), .B(n201), .C(n53), .Z(n441) );
  AOI22M1P U176 ( .A(n56), .B(\Queue[2][30] ), .C(\Queue[1][30] ), .D(n5), .Z(
        n54) );
  OAI21M1P U177 ( .A(n58), .B(n203), .C(n54), .Z(n442) );
  AOI22M1P U178 ( .A(n56), .B(\Queue[2][31] ), .C(\Queue[1][31] ), .D(n4), .Z(
        n57) );
  OAI21M1P U179 ( .A(n58), .B(n208), .C(n57), .Z(n443) );
  OAI21M1P U180 ( .A(n60), .B(n59), .C(n140), .Z(n61) );
  AOI22M1P U181 ( .A(\Queue[1][0] ), .B(n94), .C(n93), .D(Packet_Out[0]), .Z(
        n62) );
  OAI21M1P U182 ( .A(n143), .B(n8), .C(n62), .Z(n444) );
  AOI22M1P U183 ( .A(\Queue[1][1] ), .B(n94), .C(n93), .D(Packet_Out[1]), .Z(
        n63) );
  OAI21M1P U184 ( .A(n145), .B(n8), .C(n63), .Z(n445) );
  AOI22M1P U185 ( .A(\Queue[1][2] ), .B(n94), .C(n93), .D(Packet_Out[2]), .Z(
        n64) );
  OAI21M1P U186 ( .A(n147), .B(n8), .C(n64), .Z(n446) );
  AOI22M1P U187 ( .A(\Queue[1][3] ), .B(n94), .C(n93), .D(Packet_Out[3]), .Z(
        n65) );
  OAI21M1P U188 ( .A(n149), .B(n8), .C(n65), .Z(n447) );
  AOI22M1P U189 ( .A(\Queue[1][4] ), .B(n94), .C(n93), .D(Packet_Out[4]), .Z(
        n66) );
  OAI21M1P U190 ( .A(n151), .B(n8), .C(n66), .Z(n448) );
  AOI22M1P U191 ( .A(\Queue[1][5] ), .B(n94), .C(n93), .D(Packet_Out[5]), .Z(
        n67) );
  OAI21M1P U192 ( .A(n153), .B(n8), .C(n67), .Z(n449) );
  AOI22M1P U193 ( .A(\Queue[1][6] ), .B(n94), .C(n93), .D(Packet_Out[6]), .Z(
        n68) );
  OAI21M1P U194 ( .A(n155), .B(n8), .C(n68), .Z(n450) );
  AOI22M1P U195 ( .A(\Queue[1][7] ), .B(n94), .C(n93), .D(Packet_Out[7]), .Z(
        n69) );
  OAI21M1P U196 ( .A(n157), .B(n8), .C(n69), .Z(n451) );
  AOI22M1P U197 ( .A(\Queue[1][8] ), .B(n94), .C(n93), .D(Packet_Out[8]), .Z(
        n70) );
  OAI21M1P U198 ( .A(n159), .B(n8), .C(n70), .Z(n452) );
  AOI22M1P U199 ( .A(\Queue[1][9] ), .B(n94), .C(n93), .D(Packet_Out[9]), .Z(
        n71) );
  OAI21M1P U200 ( .A(n161), .B(n8), .C(n71), .Z(n453) );
  AOI22M1P U201 ( .A(\Queue[1][10] ), .B(n94), .C(n93), .D(Packet_Out[10]), 
        .Z(n72) );
  OAI21M1P U202 ( .A(n163), .B(n8), .C(n72), .Z(n454) );
  AOI22M1P U203 ( .A(\Queue[1][11] ), .B(n94), .C(n93), .D(Packet_Out[11]), 
        .Z(n73) );
  OAI21M1P U204 ( .A(n165), .B(n8), .C(n73), .Z(n455) );
  AOI22M1P U205 ( .A(\Queue[1][12] ), .B(n94), .C(n93), .D(Packet_Out[12]), 
        .Z(n74) );
  OAI21M1P U206 ( .A(n167), .B(n8), .C(n74), .Z(n456) );
  AOI22M1P U207 ( .A(\Queue[1][13] ), .B(n94), .C(n93), .D(Packet_Out[13]), 
        .Z(n75) );
  OAI21M1P U208 ( .A(n169), .B(n8), .C(n75), .Z(n457) );
  AOI22M1P U209 ( .A(\Queue[1][14] ), .B(n94), .C(n93), .D(Packet_Out[14]), 
        .Z(n76) );
  OAI21M1P U210 ( .A(n171), .B(n8), .C(n76), .Z(n458) );
  AOI22M1P U211 ( .A(\Queue[1][15] ), .B(n94), .C(n93), .D(Packet_Out[15]), 
        .Z(n77) );
  OAI21M1P U212 ( .A(n173), .B(n8), .C(n77), .Z(n459) );
  AOI22M1P U213 ( .A(\Queue[1][16] ), .B(n94), .C(n93), .D(Packet_Out[16]), 
        .Z(n78) );
  OAI21M1P U214 ( .A(n175), .B(n8), .C(n78), .Z(n460) );
  AOI22M1P U215 ( .A(\Queue[1][17] ), .B(n94), .C(n93), .D(Packet_Out[17]), 
        .Z(n79) );
  OAI21M1P U216 ( .A(n177), .B(n8), .C(n79), .Z(n461) );
  AOI22M1P U217 ( .A(\Queue[1][18] ), .B(n94), .C(n93), .D(Packet_Out[18]), 
        .Z(n80) );
  OAI21M1P U218 ( .A(n179), .B(n8), .C(n80), .Z(n462) );
  AOI22M1P U219 ( .A(\Queue[1][19] ), .B(n94), .C(n93), .D(Packet_Out[19]), 
        .Z(n81) );
  OAI21M1P U220 ( .A(n181), .B(n8), .C(n81), .Z(n463) );
  AOI22M1P U221 ( .A(\Queue[1][20] ), .B(n94), .C(n93), .D(Packet_Out[20]), 
        .Z(n82) );
  OAI21M1P U222 ( .A(n183), .B(n9), .C(n82), .Z(n464) );
  AOI22M1P U223 ( .A(\Queue[1][21] ), .B(n94), .C(n93), .D(Packet_Out[21]), 
        .Z(n83) );
  OAI21M1P U224 ( .A(n185), .B(n9), .C(n83), .Z(n465) );
  AOI22M1P U225 ( .A(\Queue[1][22] ), .B(n94), .C(n93), .D(Packet_Out[22]), 
        .Z(n84) );
  OAI21M1P U226 ( .A(n187), .B(n9), .C(n84), .Z(n466) );
  AOI22M1P U227 ( .A(\Queue[1][23] ), .B(n94), .C(n93), .D(Packet_Out[23]), 
        .Z(n85) );
  OAI21M1P U228 ( .A(n189), .B(n9), .C(n85), .Z(n467) );
  AOI22M1P U229 ( .A(\Queue[1][24] ), .B(n94), .C(n93), .D(Packet_Out[24]), 
        .Z(n86) );
  OAI21M1P U230 ( .A(n191), .B(n9), .C(n86), .Z(n468) );
  AOI22M1P U231 ( .A(\Queue[1][25] ), .B(n94), .C(n93), .D(Packet_Out[25]), 
        .Z(n87) );
  OAI21M1P U232 ( .A(n193), .B(n9), .C(n87), .Z(n469) );
  AOI22M1P U233 ( .A(\Queue[1][26] ), .B(n94), .C(n93), .D(Packet_Out[26]), 
        .Z(n88) );
  OAI21M1P U234 ( .A(n195), .B(n9), .C(n88), .Z(n470) );
  AOI22M1P U235 ( .A(\Queue[1][27] ), .B(n94), .C(n93), .D(Packet_Out[27]), 
        .Z(n89) );
  OAI21M1P U236 ( .A(n197), .B(n9), .C(n89), .Z(n471) );
  AOI22M1P U237 ( .A(\Queue[1][28] ), .B(n94), .C(n93), .D(Packet_Out[28]), 
        .Z(n90) );
  OAI21M1P U238 ( .A(n199), .B(n9), .C(n90), .Z(n472) );
  AOI22M1P U239 ( .A(\Queue[1][29] ), .B(n94), .C(n93), .D(Packet_Out[29]), 
        .Z(n91) );
  OAI21M1P U240 ( .A(n201), .B(n9), .C(n91), .Z(n473) );
  AOI22M1P U241 ( .A(\Queue[1][30] ), .B(n94), .C(n93), .D(Packet_Out[30]), 
        .Z(n92) );
  OAI21M1P U242 ( .A(n203), .B(n8), .C(n92), .Z(n474) );
  AOI22M1P U243 ( .A(\Queue[1][31] ), .B(n94), .C(n93), .D(Packet_Out[31]), 
        .Z(n95) );
  OAI21M1P U244 ( .A(n208), .B(n9), .C(n95), .Z(n475) );
  OA21M1P U245 ( .A(n138), .B(n99), .C(Rst_n), .Z(n97) );
  ND2M1P U246 ( .A(n98), .B(n136), .Z(n137) );
  AOI22M1P U247 ( .A(\Queue[2][0] ), .B(n132), .C(\Queue[3][0] ), .D(n131), 
        .Z(n100) );
  OAI21M1P U248 ( .A(n143), .B(n134), .C(n100), .Z(n476) );
  AOI22M1P U249 ( .A(\Queue[2][1] ), .B(n132), .C(n131), .D(\Queue[3][1] ), 
        .Z(n101) );
  OAI21M1P U250 ( .A(n145), .B(n134), .C(n101), .Z(n477) );
  AOI22M1P U251 ( .A(\Queue[2][2] ), .B(n132), .C(n131), .D(\Queue[3][2] ), 
        .Z(n102) );
  OAI21M1P U252 ( .A(n147), .B(n134), .C(n102), .Z(n478) );
  AOI22M1P U253 ( .A(\Queue[2][3] ), .B(n132), .C(n131), .D(\Queue[3][3] ), 
        .Z(n103) );
  OAI21M1P U254 ( .A(n149), .B(n134), .C(n103), .Z(n479) );
  AOI22M1P U255 ( .A(\Queue[2][4] ), .B(n132), .C(n131), .D(\Queue[3][4] ), 
        .Z(n104) );
  OAI21M1P U256 ( .A(n151), .B(n134), .C(n104), .Z(n480) );
  AOI22M1P U257 ( .A(\Queue[2][5] ), .B(n132), .C(n131), .D(\Queue[3][5] ), 
        .Z(n105) );
  OAI21M1P U258 ( .A(n153), .B(n134), .C(n105), .Z(n481) );
  AOI22M1P U259 ( .A(\Queue[2][6] ), .B(n132), .C(n131), .D(\Queue[3][6] ), 
        .Z(n106) );
  OAI21M1P U260 ( .A(n155), .B(n134), .C(n106), .Z(n482) );
  AOI22M1P U261 ( .A(\Queue[2][7] ), .B(n132), .C(n131), .D(\Queue[3][7] ), 
        .Z(n107) );
  OAI21M1P U262 ( .A(n157), .B(n134), .C(n107), .Z(n483) );
  AOI22M1P U263 ( .A(\Queue[2][8] ), .B(n132), .C(n131), .D(\Queue[3][8] ), 
        .Z(n108) );
  OAI21M1P U264 ( .A(n159), .B(n134), .C(n108), .Z(n484) );
  AOI22M1P U265 ( .A(\Queue[2][9] ), .B(n132), .C(n131), .D(\Queue[3][9] ), 
        .Z(n109) );
  OAI21M1P U266 ( .A(n161), .B(n134), .C(n109), .Z(n485) );
  AOI22M1P U267 ( .A(\Queue[2][10] ), .B(n132), .C(n131), .D(\Queue[3][10] ), 
        .Z(n110) );
  OAI21M1P U268 ( .A(n163), .B(n134), .C(n110), .Z(n486) );
  AOI22M1P U269 ( .A(\Queue[2][11] ), .B(n132), .C(n131), .D(\Queue[3][11] ), 
        .Z(n111) );
  OAI21M1P U270 ( .A(n165), .B(n134), .C(n111), .Z(n487) );
  AOI22M1P U271 ( .A(\Queue[2][12] ), .B(n132), .C(n131), .D(\Queue[3][12] ), 
        .Z(n112) );
  OAI21M1P U272 ( .A(n167), .B(n134), .C(n112), .Z(n488) );
  AOI22M1P U273 ( .A(\Queue[2][13] ), .B(n132), .C(n131), .D(\Queue[3][13] ), 
        .Z(n113) );
  OAI21M1P U274 ( .A(n169), .B(n134), .C(n113), .Z(n489) );
  AOI22M1P U275 ( .A(\Queue[2][14] ), .B(n132), .C(n131), .D(\Queue[3][14] ), 
        .Z(n114) );
  OAI21M1P U276 ( .A(n171), .B(n134), .C(n114), .Z(n490) );
  AOI22M1P U277 ( .A(\Queue[2][15] ), .B(n132), .C(n131), .D(\Queue[3][15] ), 
        .Z(n115) );
  OAI21M1P U278 ( .A(n173), .B(n134), .C(n115), .Z(n491) );
  AOI22M1P U279 ( .A(\Queue[2][16] ), .B(n132), .C(n131), .D(\Queue[3][16] ), 
        .Z(n116) );
  OAI21M1P U280 ( .A(n175), .B(n134), .C(n116), .Z(n492) );
  AOI22M1P U281 ( .A(\Queue[2][17] ), .B(n132), .C(n131), .D(\Queue[3][17] ), 
        .Z(n117) );
  OAI21M1P U282 ( .A(n177), .B(n134), .C(n117), .Z(n493) );
  AOI22M1P U283 ( .A(\Queue[2][18] ), .B(n132), .C(n131), .D(\Queue[3][18] ), 
        .Z(n118) );
  OAI21M1P U284 ( .A(n179), .B(n134), .C(n118), .Z(n494) );
  AOI22M1P U285 ( .A(\Queue[2][19] ), .B(n132), .C(n131), .D(\Queue[3][19] ), 
        .Z(n119) );
  OAI21M1P U286 ( .A(n181), .B(n134), .C(n119), .Z(n495) );
  AOI22M1P U287 ( .A(\Queue[2][20] ), .B(n132), .C(n131), .D(\Queue[3][20] ), 
        .Z(n120) );
  OAI21M1P U288 ( .A(n183), .B(n134), .C(n120), .Z(n496) );
  AOI22M1P U289 ( .A(\Queue[2][21] ), .B(n132), .C(n131), .D(\Queue[3][21] ), 
        .Z(n121) );
  OAI21M1P U290 ( .A(n185), .B(n134), .C(n121), .Z(n497) );
  AOI22M1P U291 ( .A(\Queue[2][22] ), .B(n132), .C(n131), .D(\Queue[3][22] ), 
        .Z(n122) );
  OAI21M1P U292 ( .A(n187), .B(n134), .C(n122), .Z(n498) );
  AOI22M1P U293 ( .A(\Queue[2][23] ), .B(n132), .C(n131), .D(\Queue[3][23] ), 
        .Z(n123) );
  OAI21M1P U294 ( .A(n189), .B(n134), .C(n123), .Z(n499) );
  AOI22M1P U295 ( .A(\Queue[2][24] ), .B(n132), .C(n131), .D(\Queue[3][24] ), 
        .Z(n124) );
  OAI21M1P U296 ( .A(n191), .B(n134), .C(n124), .Z(n500) );
  AOI22M1P U297 ( .A(\Queue[2][25] ), .B(n132), .C(n131), .D(\Queue[3][25] ), 
        .Z(n125) );
  OAI21M1P U298 ( .A(n193), .B(n134), .C(n125), .Z(n501) );
  AOI22M1P U299 ( .A(\Queue[2][26] ), .B(n132), .C(n131), .D(\Queue[3][26] ), 
        .Z(n126) );
  OAI21M1P U300 ( .A(n195), .B(n134), .C(n126), .Z(n502) );
  AOI22M1P U301 ( .A(\Queue[2][27] ), .B(n132), .C(n131), .D(\Queue[3][27] ), 
        .Z(n127) );
  OAI21M1P U302 ( .A(n197), .B(n134), .C(n127), .Z(n503) );
  AOI22M1P U303 ( .A(\Queue[2][28] ), .B(n132), .C(n131), .D(\Queue[3][28] ), 
        .Z(n128) );
  OAI21M1P U304 ( .A(n199), .B(n134), .C(n128), .Z(n504) );
  AOI22M1P U305 ( .A(\Queue[2][29] ), .B(n132), .C(n131), .D(\Queue[3][29] ), 
        .Z(n129) );
  OAI21M1P U306 ( .A(n201), .B(n134), .C(n129), .Z(n505) );
  AOI22M1P U307 ( .A(\Queue[2][30] ), .B(n132), .C(n131), .D(\Queue[3][30] ), 
        .Z(n130) );
  OAI21M1P U308 ( .A(n203), .B(n134), .C(n130), .Z(n506) );
  AOI22M1P U309 ( .A(\Queue[2][31] ), .B(n132), .C(n131), .D(\Queue[3][31] ), 
        .Z(n133) );
  OAI21M1P U310 ( .A(n208), .B(n134), .C(n133), .Z(n507) );
  OA21M1P U311 ( .A(n138), .B(n139), .C(Rst_n), .Z(n135) );
  AOI22M1P U312 ( .A(\Queue[3][0] ), .B(n10), .C(n204), .D(\Queue[4][0] ), .Z(
        n142) );
  OAI21M1P U313 ( .A(n143), .B(n207), .C(n142), .Z(n508) );
  AOI22M1P U314 ( .A(\Queue[3][1] ), .B(n10), .C(n204), .D(\Queue[4][1] ), .Z(
        n144) );
  OAI21M1P U315 ( .A(n145), .B(n207), .C(n144), .Z(n509) );
  AOI22M1P U316 ( .A(\Queue[3][2] ), .B(n10), .C(n204), .D(\Queue[4][2] ), .Z(
        n146) );
  OAI21M1P U317 ( .A(n147), .B(n207), .C(n146), .Z(n510) );
  AOI22M1P U318 ( .A(\Queue[3][3] ), .B(n10), .C(n204), .D(\Queue[4][3] ), .Z(
        n148) );
  OAI21M1P U319 ( .A(n149), .B(n207), .C(n148), .Z(n511) );
  AOI22M1P U320 ( .A(\Queue[3][4] ), .B(n10), .C(n204), .D(\Queue[4][4] ), .Z(
        n150) );
  OAI21M1P U321 ( .A(n151), .B(n207), .C(n150), .Z(n512) );
  AOI22M1P U322 ( .A(\Queue[3][5] ), .B(n10), .C(n204), .D(\Queue[4][5] ), .Z(
        n152) );
  OAI21M1P U323 ( .A(n153), .B(n207), .C(n152), .Z(n513) );
  AOI22M1P U324 ( .A(\Queue[3][6] ), .B(n10), .C(n204), .D(\Queue[4][6] ), .Z(
        n154) );
  OAI21M1P U325 ( .A(n155), .B(n207), .C(n154), .Z(n514) );
  AOI22M1P U326 ( .A(\Queue[3][7] ), .B(n10), .C(n204), .D(\Queue[4][7] ), .Z(
        n156) );
  OAI21M1P U327 ( .A(n157), .B(n207), .C(n156), .Z(n515) );
  AOI22M1P U328 ( .A(\Queue[3][8] ), .B(n10), .C(n204), .D(\Queue[4][8] ), .Z(
        n158) );
  OAI21M1P U329 ( .A(n159), .B(n207), .C(n158), .Z(n516) );
  AOI22M1P U330 ( .A(\Queue[3][9] ), .B(n10), .C(n204), .D(\Queue[4][9] ), .Z(
        n160) );
  OAI21M1P U331 ( .A(n161), .B(n207), .C(n160), .Z(n517) );
  AOI22M1P U332 ( .A(\Queue[3][10] ), .B(n10), .C(n204), .D(\Queue[4][10] ), 
        .Z(n162) );
  OAI21M1P U333 ( .A(n163), .B(n207), .C(n162), .Z(n518) );
  AOI22M1P U334 ( .A(\Queue[3][11] ), .B(n10), .C(n204), .D(\Queue[4][11] ), 
        .Z(n164) );
  OAI21M1P U335 ( .A(n165), .B(n207), .C(n164), .Z(n519) );
  AOI22M1P U336 ( .A(\Queue[3][12] ), .B(n10), .C(n204), .D(\Queue[4][12] ), 
        .Z(n166) );
  OAI21M1P U337 ( .A(n167), .B(n207), .C(n166), .Z(n520) );
  AOI22M1P U338 ( .A(\Queue[3][13] ), .B(n10), .C(n204), .D(\Queue[4][13] ), 
        .Z(n168) );
  OAI21M1P U339 ( .A(n169), .B(n207), .C(n168), .Z(n521) );
  AOI22M1P U340 ( .A(\Queue[3][14] ), .B(n10), .C(n204), .D(\Queue[4][14] ), 
        .Z(n170) );
  OAI21M1P U341 ( .A(n171), .B(n207), .C(n170), .Z(n522) );
  AOI22M1P U342 ( .A(\Queue[3][15] ), .B(n10), .C(n204), .D(\Queue[4][15] ), 
        .Z(n172) );
  OAI21M1P U343 ( .A(n173), .B(n207), .C(n172), .Z(n523) );
  AOI22M1P U344 ( .A(\Queue[3][16] ), .B(n10), .C(n204), .D(\Queue[4][16] ), 
        .Z(n174) );
  OAI21M1P U345 ( .A(n175), .B(n207), .C(n174), .Z(n524) );
  AOI22M1P U346 ( .A(\Queue[3][17] ), .B(n10), .C(n204), .D(\Queue[4][17] ), 
        .Z(n176) );
  OAI21M1P U347 ( .A(n177), .B(n207), .C(n176), .Z(n525) );
  AOI22M1P U348 ( .A(\Queue[3][18] ), .B(n10), .C(n204), .D(\Queue[4][18] ), 
        .Z(n178) );
  OAI21M1P U349 ( .A(n179), .B(n207), .C(n178), .Z(n526) );
  AOI22M1P U350 ( .A(\Queue[3][19] ), .B(n10), .C(n204), .D(\Queue[4][19] ), 
        .Z(n180) );
  OAI21M1P U351 ( .A(n181), .B(n207), .C(n180), .Z(n527) );
  AOI22M1P U352 ( .A(\Queue[3][20] ), .B(n11), .C(n204), .D(\Queue[4][20] ), 
        .Z(n182) );
  OAI21M1P U353 ( .A(n183), .B(n207), .C(n182), .Z(n528) );
  AOI22M1P U354 ( .A(\Queue[3][21] ), .B(n11), .C(n204), .D(\Queue[4][21] ), 
        .Z(n184) );
  OAI21M1P U355 ( .A(n185), .B(n207), .C(n184), .Z(n529) );
  AOI22M1P U356 ( .A(\Queue[3][22] ), .B(n11), .C(n204), .D(\Queue[4][22] ), 
        .Z(n186) );
  OAI21M1P U357 ( .A(n187), .B(n207), .C(n186), .Z(n530) );
  AOI22M1P U358 ( .A(\Queue[3][23] ), .B(n11), .C(n204), .D(\Queue[4][23] ), 
        .Z(n188) );
  OAI21M1P U359 ( .A(n189), .B(n207), .C(n188), .Z(n531) );
  AOI22M1P U360 ( .A(\Queue[3][24] ), .B(n11), .C(n204), .D(\Queue[4][24] ), 
        .Z(n190) );
  OAI21M1P U361 ( .A(n191), .B(n207), .C(n190), .Z(n532) );
  AOI22M1P U362 ( .A(\Queue[3][25] ), .B(n11), .C(n204), .D(\Queue[4][25] ), 
        .Z(n192) );
  OAI21M1P U363 ( .A(n193), .B(n207), .C(n192), .Z(n533) );
  AOI22M1P U364 ( .A(\Queue[3][26] ), .B(n11), .C(n204), .D(\Queue[4][26] ), 
        .Z(n194) );
  OAI21M1P U365 ( .A(n195), .B(n207), .C(n194), .Z(n534) );
  AOI22M1P U366 ( .A(\Queue[3][27] ), .B(n11), .C(n204), .D(\Queue[4][27] ), 
        .Z(n196) );
  OAI21M1P U367 ( .A(n197), .B(n207), .C(n196), .Z(n535) );
  AOI22M1P U368 ( .A(\Queue[3][28] ), .B(n11), .C(n204), .D(\Queue[4][28] ), 
        .Z(n198) );
  OAI21M1P U369 ( .A(n199), .B(n207), .C(n198), .Z(n536) );
  AOI22M1P U370 ( .A(\Queue[3][29] ), .B(n11), .C(n204), .D(\Queue[4][29] ), 
        .Z(n200) );
  OAI21M1P U371 ( .A(n201), .B(n207), .C(n200), .Z(n537) );
  AOI22M1P U372 ( .A(\Queue[3][30] ), .B(n10), .C(n204), .D(\Queue[4][30] ), 
        .Z(n202) );
  OAI21M1P U373 ( .A(n203), .B(n207), .C(n202), .Z(n538) );
  AOI22M1P U374 ( .A(\Queue[3][31] ), .B(n11), .C(n204), .D(\Queue[4][31] ), 
        .Z(n206) );
  OAI21M1P U375 ( .A(n208), .B(n207), .C(n206), .Z(n539) );
  N1M1P U376 ( .A(n540), .Z(Empty) );
  AOI22M1P U377 ( .A(n375), .B(n374), .C(n373), .D(Empty), .Z(n541) );
endmodule


module Link_Control_3 ( Clk_r, Rst_n, Tx_Ready, Tx_Error, RxData_Valid, RxData, 
        Packet_From_Core, TxQueue_Write, RxQueue_Read, TxData_Valid, TxData, 
        Error_Ack, Core_Rcv_Ready, Packet_To_Core, RxQueue_Empty, TxQueue_Full
 );
  input [31:0] RxData;
  input [31:0] Packet_From_Core;
  output [31:0] TxData;
  output [31:0] Packet_To_Core;
  input Clk_r, Rst_n, Tx_Ready, Tx_Error, RxData_Valid, TxQueue_Write,
         RxQueue_Read;
  output TxData_Valid, Error_Ack, Core_Rcv_Ready, RxQueue_Empty, TxQueue_Full;
  wire   TxQueue_Read, TxQueue_Empty, RxQueue_Write, RxQueue_Full, N9, N16, n5,
         n6, n7, n8, n9;

  Packet_Queue_8 TxQueue ( .Clk_r(Clk_r), .Rst_n(Rst_n), .Packet_In(
        Packet_From_Core), .Read_Ack(TxQueue_Read), .Write_Ack(TxQueue_Write), 
        .Packet_Out(TxData), .Empty(TxQueue_Empty), .Full(TxQueue_Full) );
  Packet_Queue_7 RxQueue ( .Clk_r(Clk_r), .Rst_n(Rst_n), .Packet_In(RxData), 
        .Read_Ack(RxQueue_Read), .Write_Ack(RxQueue_Write), .Packet_Out(
        Packet_To_Core), .Empty(RxQueue_Empty), .Full(RxQueue_Full) );
  FD2QM1P Core_Rcv_Ready_reg ( .D(N9), .CP(Clk_r), .CD(Rst_n), .Q(
        Core_Rcv_Ready) );
  FD2QM1P TxQueue_Read_reg ( .D(N16), .CP(Clk_r), .CD(Rst_n), .Q(TxQueue_Read)
         );
  FD4QM1P RxQueue_Write_reg ( .D(n7), .CP(Clk_r), .SD(Rst_n), .Q(n6) );
  FD4QM1P TxData_Valid_reg ( .D(n9), .CP(Clk_r), .SD(Rst_n), .Q(n8) );
  N1M3P U3 ( .A(n6), .Z(RxQueue_Write) );
  NR2M1P U4 ( .A(n8), .B(Tx_Ready), .Z(N16) );
  NR2M1P U5 ( .A(RxData_Valid), .B(RxQueue_Full), .Z(n5) );
  OA21M1P U6 ( .A(Core_Rcv_Ready), .B(n5), .C(n6), .Z(N9) );
  N1M1P U7 ( .A(n8), .Z(TxData_Valid) );
  ND3M1P U8 ( .A(n6), .B(Core_Rcv_Ready), .C(RxData_Valid), .Z(n7) );
  AO21CNM1P U9 ( .A(n8), .B(TxQueue_Empty), .C(Tx_Ready), .Z(n9) );
endmodule


module core ( Clk_r, Rst_n, N_Tx_Ready, N_Tx_Error, N_RxData_Valid, N_RxData, 
        S_Tx_Ready, S_Tx_Error, S_RxData_Valid, S_RxData, W_Tx_Ready, 
        W_Tx_Error, W_RxData_Valid, W_RxData, E_Tx_Ready, E_Tx_Error, 
        E_RxData_Valid, E_RxData, Packet_From_Node, Packet_From_Node_Valid, 
        N_TxData_Valid, N_TxData, N_Error_Ack, N_Core_Rcv_Ready, 
        S_TxData_Valid, S_TxData, S_Error_Ack, S_Core_Rcv_Ready, 
        W_TxData_Valid, W_TxData, W_Error_Ack, W_Core_Rcv_Ready, 
        E_TxData_Valid, E_TxData, E_Error_Ack, E_Core_Rcv_Ready, Core_Load_Ack, 
        Packet_To_Node, Packet_To_Node_Valid );
  input [31:0] N_RxData;
  input [31:0] S_RxData;
  input [31:0] W_RxData;
  input [31:0] E_RxData;
  input [31:0] Packet_From_Node;
  output [31:0] N_TxData;
  output [31:0] S_TxData;
  output [31:0] W_TxData;
  output [31:0] E_TxData;
  output [31:0] Packet_To_Node;
  input Clk_r, Rst_n, N_Tx_Ready, N_Tx_Error, N_RxData_Valid, S_Tx_Ready,
         S_Tx_Error, S_RxData_Valid, W_Tx_Ready, W_Tx_Error, W_RxData_Valid,
         E_Tx_Ready, E_Tx_Error, E_RxData_Valid, Packet_From_Node_Valid;
  output N_TxData_Valid, N_Error_Ack, N_Core_Rcv_Ready, S_TxData_Valid,
         S_Error_Ack, S_Core_Rcv_Ready, W_TxData_Valid, W_Error_Ack,
         W_Core_Rcv_Ready, E_TxData_Valid, E_Error_Ack, E_Core_Rcv_Ready,
         Core_Load_Ack, Packet_To_Node_Valid;
  wire   N_TxQueue_Write, N_RxQueue_Read, N_RxQueue_Empty, N_TxQueue_Full,
         S_TxQueue_Write, S_RxQueue_Read, S_RxQueue_Empty, S_TxQueue_Full,
         E_TxQueue_Write, E_RxQueue_Read, E_RxQueue_Empty, E_TxQueue_Full,
         W_TxQueue_Write, W_RxQueue_Read, W_RxQueue_Empty, W_TxQueue_Full,
         NM_Empty, NM_Full, NM_Read, NM_Write;
  wire   [31:0] N_Tx_Packet;
  wire   [31:0] N_Rx_Packet;
  wire   [31:0] S_Tx_Packet;
  wire   [31:0] S_Rx_Packet;
  wire   [31:0] E_Tx_Packet;
  wire   [31:0] E_Rx_Packet;
  wire   [31:0] W_Tx_Packet;
  wire   [31:0] W_Rx_Packet;
  wire   [7:0] Router_Addr;
  wire   [3:0] Link_Config;
  wire   [31:0] NM_In_Packet;
  wire   [31:0] NM_Out_Packet;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7;

  Link_Control_0 N_Link_Control ( .Clk_r(Clk_r), .Rst_n(Rst_n), .Tx_Ready(
        N_Tx_Ready), .Tx_Error(1'b0), .RxData_Valid(N_RxData_Valid), .RxData(
        N_RxData), .Packet_From_Core(N_Tx_Packet), .TxQueue_Write(
        N_TxQueue_Write), .RxQueue_Read(N_RxQueue_Read), .TxData_Valid(
        N_TxData_Valid), .TxData(N_TxData), .Core_Rcv_Ready(N_Core_Rcv_Ready), 
        .Packet_To_Core(N_Rx_Packet), .RxQueue_Empty(N_RxQueue_Empty), 
        .TxQueue_Full(N_TxQueue_Full) );
  Link_Control_3 S_Link_Control ( .Clk_r(Clk_r), .Rst_n(Rst_n), .Tx_Ready(
        S_Tx_Ready), .Tx_Error(1'b0), .RxData_Valid(S_RxData_Valid), .RxData(
        S_RxData), .Packet_From_Core(S_Tx_Packet), .TxQueue_Write(
        S_TxQueue_Write), .RxQueue_Read(S_RxQueue_Read), .TxData_Valid(
        S_TxData_Valid), .TxData(S_TxData), .Core_Rcv_Ready(S_Core_Rcv_Ready), 
        .Packet_To_Core(S_Rx_Packet), .RxQueue_Empty(S_RxQueue_Empty), 
        .TxQueue_Full(S_TxQueue_Full) );
  Link_Control_2 E_Link_Control ( .Clk_r(Clk_r), .Rst_n(Rst_n), .Tx_Ready(
        E_Tx_Ready), .Tx_Error(1'b0), .RxData_Valid(E_RxData_Valid), .RxData(
        E_RxData), .Packet_From_Core(E_Tx_Packet), .TxQueue_Write(
        E_TxQueue_Write), .RxQueue_Read(E_RxQueue_Read), .TxData_Valid(
        E_TxData_Valid), .TxData(E_TxData), .Core_Rcv_Ready(E_Core_Rcv_Ready), 
        .Packet_To_Core(E_Rx_Packet), .RxQueue_Empty(E_RxQueue_Empty), 
        .TxQueue_Full(E_TxQueue_Full) );
  Link_Control_1 W_Link_Control ( .Clk_r(Clk_r), .Rst_n(Rst_n), .Tx_Ready(
        W_Tx_Ready), .Tx_Error(1'b0), .RxData_Valid(W_RxData_Valid), .RxData(
        W_RxData), .Packet_From_Core(W_Tx_Packet), .TxQueue_Write(
        W_TxQueue_Write), .RxQueue_Read(W_RxQueue_Read), .TxData_Valid(
        W_TxData_Valid), .TxData(W_TxData), .Core_Rcv_Ready(W_Core_Rcv_Ready), 
        .Packet_To_Core(W_Rx_Packet), .RxQueue_Empty(W_RxQueue_Empty), 
        .TxQueue_Full(W_TxQueue_Full) );
  Routing_State_Machine routing_state_machine ( .Clk_r(Clk_r), .Rst_n(Rst_n), 
        .Router_Address(Router_Addr), .Link_Config(Link_Config), 
        .Packet_From_Link_N(N_Rx_Packet), .Packet_From_Link_S(S_Rx_Packet), 
        .Packet_From_Link_W(W_Rx_Packet), .Packet_From_Link_E(E_Rx_Packet), 
        .Packet_From_Node({NM_In_Packet[31:24], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, NM_In_Packet[15:0]}), .RxQueue_Empty_N(
        N_RxQueue_Empty), .RxQueue_Empty_S(S_RxQueue_Empty), .RxQueue_Empty_W(
        W_RxQueue_Empty), .RxQueue_Empty_E(E_RxQueue_Empty), .TxQueue_Full_N(
        N_TxQueue_Full), .TxQueue_Full_S(S_TxQueue_Full), .TxQueue_Full_W(
        W_TxQueue_Full), .TxQueue_Full_E(E_TxQueue_Full), .To_Node_Full(
        NM_Full), .Node_Queue_Empty(NM_Empty), .Packet_To_Link_N(N_Tx_Packet), 
        .Packet_To_Link_S(S_Tx_Packet), .Packet_To_Link_W(W_Tx_Packet), 
        .Packet_To_Link_E(E_Tx_Packet), .Packet_To_Node(NM_Out_Packet), 
        .TxQueue_Write_N(N_TxQueue_Write), .TxQueue_Write_S(S_TxQueue_Write), 
        .TxQueue_Write_W(W_TxQueue_Write), .TxQueue_Write_E(E_TxQueue_Write), 
        .To_Node_Write(NM_Write), .RxQueue_Read_N(N_RxQueue_Read), 
        .RxQueue_Read_S(S_RxQueue_Read), .RxQueue_Read_W(W_RxQueue_Read), 
        .RxQueue_Read_E(E_RxQueue_Read), .Node_Read(NM_Read) );
  Node_Manager node_manager ( .Clk_r(Clk_r), .Rst_n(Rst_n), .Packet_From_Core(
        NM_Out_Packet), .Packet_From_Node(Packet_From_Node), 
        .Packet_From_Node_Valid(Packet_From_Node_Valid), .Read_Packet(NM_Read), 
        .To_Node_Write(NM_Write), .Router_Address(Router_Addr), .Link_Config(
        Link_Config), .Packet_To_Core({NM_In_Packet[31:24], 
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, NM_In_Packet[15:0]}), 
        .Packet_To_Node(Packet_To_Node), .Packet_To_Node_Valid(
        Packet_To_Node_Valid), .Core_Load_Ack(Core_Load_Ack), .Queue_Empty(
        NM_Empty), .To_Node_Full(NM_Full) );
endmodule


module tx_0 ( Clk_s, Rst_n, TxData_Valid, TxData, Error_Ack, Rx_Ready, 
        Rx_Error, Tx_Ready, Tx_Error, S_Data );
  input [31:0] TxData;
  input Clk_s, Rst_n, TxData_Valid, Error_Ack, Rx_Ready, Rx_Error;
  output Tx_Ready, Tx_Error, S_Data;
  wire   N100, N101, N102, N103, N104, N105, N106, N107, N108, N109, N110,
         N111, N112, N113, N114, N115, N116, N117, N118, N119, N120, N121,
         N122, N123, N124, N125, N126, N127, N128, N129, N130, N131, N132,
         N146, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n23, n24, n25, n26, n27, n28, n93, n157, n162, n17, n18,
         n19, n20, n21, n22, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142;
  wire   [32:0] transmissionPacket;
  wire   [5:0] bitCount;

  FD4QM1P zeroPatternDetected_reg ( .D(n14), .CP(Clk_s), .SD(Rst_n), .Q(n15)
         );
  FD4QM1P DataTxInProg_reg ( .D(n12), .CP(Clk_s), .SD(Rst_n), .Q(n13) );
  FD4QM1P Tx_Ready_reg ( .D(n162), .CP(Clk_s), .SD(Rst_n), .Q(Tx_Ready) );
  FD2LQM1P \transmissionPacket_reg[1]  ( .D(TxData[0]), .LD(n58), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[1]) );
  FD2LQM1P \transmissionPacket_reg[2]  ( .D(TxData[1]), .LD(n58), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[2]) );
  FD2LQM1P \transmissionPacket_reg[3]  ( .D(TxData[2]), .LD(n58), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[3]) );
  FD2LQM1P \transmissionPacket_reg[4]  ( .D(TxData[3]), .LD(n58), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[4]) );
  FD2LQM1P \transmissionPacket_reg[5]  ( .D(TxData[4]), .LD(n58), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[5]) );
  FD2LQM1P \transmissionPacket_reg[6]  ( .D(TxData[5]), .LD(n58), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[6]) );
  FD2LQM1P \transmissionPacket_reg[7]  ( .D(TxData[6]), .LD(n58), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[7]) );
  FD2LQM1P \transmissionPacket_reg[8]  ( .D(TxData[7]), .LD(n58), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[8]) );
  FD2LQM1P \transmissionPacket_reg[9]  ( .D(TxData[8]), .LD(n58), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[9]) );
  FD2LQM1P \transmissionPacket_reg[10]  ( .D(TxData[9]), .LD(n58), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[10]) );
  FD2LQM1P \transmissionPacket_reg[11]  ( .D(TxData[10]), .LD(n58), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[11]) );
  FD2LQM1P \transmissionPacket_reg[12]  ( .D(TxData[11]), .LD(n58), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[12]) );
  FD2LQM1P \transmissionPacket_reg[13]  ( .D(TxData[12]), .LD(n58), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[13]) );
  FD2LQM1P \transmissionPacket_reg[14]  ( .D(TxData[13]), .LD(n58), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[14]) );
  FD2LQM1P \transmissionPacket_reg[15]  ( .D(TxData[14]), .LD(n58), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[15]) );
  FD2LQM1P \transmissionPacket_reg[16]  ( .D(TxData[15]), .LD(n58), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[16]) );
  FD2LQM1P \transmissionPacket_reg[17]  ( .D(TxData[16]), .LD(n58), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[17]) );
  FD2LQM1P \transmissionPacket_reg[18]  ( .D(TxData[17]), .LD(n58), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[18]) );
  FD2LQM1P \transmissionPacket_reg[19]  ( .D(TxData[18]), .LD(n58), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[19]) );
  FD2LQM1P \transmissionPacket_reg[20]  ( .D(TxData[19]), .LD(n58), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[20]) );
  FD2LQM1P \transmissionPacket_reg[21]  ( .D(TxData[20]), .LD(n58), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[21]) );
  FD2LQM1P \transmissionPacket_reg[22]  ( .D(TxData[21]), .LD(n58), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[22]) );
  FD2LQM1P \transmissionPacket_reg[23]  ( .D(TxData[22]), .LD(n16), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[23]) );
  FD2LQM1P \transmissionPacket_reg[24]  ( .D(TxData[23]), .LD(n16), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[24]) );
  FD2LQM1P \transmissionPacket_reg[25]  ( .D(TxData[24]), .LD(n16), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[25]) );
  FD2LQM1P \transmissionPacket_reg[26]  ( .D(TxData[25]), .LD(n16), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[26]) );
  FD2LQM1P \transmissionPacket_reg[27]  ( .D(TxData[26]), .LD(n16), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[27]) );
  FD2LQM1P \transmissionPacket_reg[28]  ( .D(TxData[27]), .LD(n16), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[28]) );
  FD2LQM1P \transmissionPacket_reg[29]  ( .D(TxData[28]), .LD(n16), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[29]) );
  FD2LQM1P \transmissionPacket_reg[30]  ( .D(TxData[29]), .LD(n16), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[30]) );
  FD2LQM1P \transmissionPacket_reg[31]  ( .D(TxData[30]), .LD(n16), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[31]) );
  FD2LQM1P \transmissionPacket_reg[32]  ( .D(TxData[31]), .LD(n58), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[32]) );
  FD4QM1P \startSequenceCount_reg[1]  ( .D(n10), .CP(Clk_s), .SD(Rst_n), .Q(
        n11) );
  FD4QM1P \startSequenceCount_reg[2]  ( .D(n8), .CP(Clk_s), .SD(Rst_n), .Q(n9)
         );
  FD4QM1P \startSequenceCount_reg[0]  ( .D(n6), .CP(Clk_s), .SD(Rst_n), .Q(n7)
         );
  FD4QM1P startSequence_reg ( .D(n93), .CP(Clk_s), .SD(Rst_n), .Q(n5) );
  FD4QM1P \zeroCount_reg[0]  ( .D(n3), .CP(Clk_s), .SD(Rst_n), .Q(n4) );
  FD4QM1P \zeroCount_reg[1]  ( .D(n1), .CP(Clk_s), .SD(Rst_n), .Q(n2) );
  FD4QM1P S_Data_reg ( .D(N146), .CP(Clk_s), .SD(Rst_n), .Q(S_Data) );
  FD2QM1P \bitCount_reg[0]  ( .D(n23), .CP(Clk_s), .CD(Rst_n), .Q(bitCount[0])
         );
  FD2QM1P \bitCount_reg[3]  ( .D(n26), .CP(Clk_s), .CD(Rst_n), .Q(bitCount[3])
         );
  FD2QM1P \bitCount_reg[1]  ( .D(n24), .CP(Clk_s), .CD(Rst_n), .Q(bitCount[1])
         );
  FD2QM1P \bitCount_reg[4]  ( .D(n27), .CP(Clk_s), .CD(Rst_n), .Q(bitCount[4])
         );
  FD2QM1P \bitCount_reg[5]  ( .D(n28), .CP(Clk_s), .CD(Rst_n), .Q(bitCount[5])
         );
  FD2QM1P \bitCount_reg[2]  ( .D(n25), .CP(Clk_s), .CD(Rst_n), .Q(bitCount[2])
         );
  FD2QM1P \transmissionPacket_reg[0]  ( .D(n157), .CP(Clk_s), .CD(Rst_n), .Q(
        transmissionPacket[0]) );
  NR2BNM1P U3 ( .B(bitCount[4]), .A(bitCount[5]), .Z(n46) );
  ND2BNM1P U4 ( .B(bitCount[1]), .A(bitCount[0]), .Z(n55) );
  ND2BNM1P U5 ( .B(bitCount[0]), .A(bitCount[1]), .Z(n18) );
  N1M1P U6 ( .A(bitCount[2]), .Z(n124) );
  ND4M1P U7 ( .A(n15), .B(n5), .C(n138), .D(n81), .Z(n131) );
  AND2M1P U8 ( .A(Tx_Ready), .B(TxData_Valid), .Z(n16) );
  AOI22DNM1P U9 ( .A(n2), .B(n142), .D(n140), .C(n141), .Z(n17) );
  OA21M1P U10 ( .A(n2), .B(n20), .C(n17), .Z(n1) );
  N1M1P U11 ( .A(n131), .Z(n133) );
  NR3M1P U12 ( .A(n37), .B(n36), .C(n35), .Z(n40) );
  OR2M1P U13 ( .A(bitCount[0]), .B(bitCount[1]), .Z(n54) );
  BUFM2P U14 ( .A(n16), .Z(n58) );
  ND2BNM1P U15 ( .B(n19), .A(n4), .Z(n20) );
  NR2M1P U16 ( .A(n19), .B(n4), .Z(n142) );
  N1M1P U17 ( .A(bitCount[3]), .Z(n57) );
  ND2M1P U18 ( .A(n48), .B(n46), .Z(n43) );
  OA21M1P U19 ( .A(n4), .B(n140), .C(n20), .Z(n3) );
  NR2M1P U20 ( .A(n18), .B(n52), .Z(N106) );
  NR2M1P U21 ( .A(n18), .B(n47), .Z(N130) );
  NR2M1P U22 ( .A(n50), .B(n18), .Z(N102) );
  NR2M1P U23 ( .A(n18), .B(n45), .Z(N126) );
  NR2M1P U24 ( .A(n18), .B(n44), .Z(N122) );
  NR2M1P U25 ( .A(n18), .B(n43), .Z(N118) );
  NR2M1P U26 ( .A(n18), .B(n42), .Z(N114) );
  NR2M1P U27 ( .A(n56), .B(n18), .Z(N110) );
  ND2M1P U28 ( .A(n41), .B(n40), .Z(n19) );
  AOI22M1P U29 ( .A(transmissionPacket[13]), .B(N119), .C(
        transmissionPacket[12]), .D(N120), .Z(n21) );
  AOI22M1P U30 ( .A(transmissionPacket[22]), .B(N110), .C(
        transmissionPacket[21]), .D(N111), .Z(n22) );
  AOI22M1P U31 ( .A(transmissionPacket[23]), .B(N109), .C(
        transmissionPacket[20]), .D(N112), .Z(n29) );
  AOI22M1P U32 ( .A(transmissionPacket[2]), .B(N130), .C(transmissionPacket[1]), .D(N131), .Z(n30) );
  AOI22M1P U33 ( .A(transmissionPacket[4]), .B(N128), .C(transmissionPacket[6]), .D(N126), .Z(n31) );
  AOI22M1P U34 ( .A(transmissionPacket[5]), .B(N127), .C(transmissionPacket[3]), .D(N129), .Z(n32) );
  AOI22M1P U35 ( .A(transmissionPacket[7]), .B(N125), .C(transmissionPacket[9]), .D(N123), .Z(n33) );
  AOI22M1P U36 ( .A(transmissionPacket[11]), .B(N121), .C(
        transmissionPacket[10]), .D(N122), .Z(n34) );
  ND4M1P U37 ( .A(n69), .B(n68), .C(n67), .D(n21), .Z(n35) );
  ND4M1P U38 ( .A(n65), .B(n64), .C(n29), .D(n22), .Z(n36) );
  ND4M1P U39 ( .A(n30), .B(n60), .C(n59), .D(n66), .Z(n37) );
  ND4M1P U40 ( .A(n34), .B(n33), .C(n32), .D(n31), .Z(n38) );
  ND3M1P U41 ( .A(n138), .B(n15), .C(n5), .Z(n39) );
  AOI211M1P U42 ( .A(N124), .B(transmissionPacket[8]), .C(n39), .D(n38), .Z(
        n41) );
  NR2M1P U43 ( .A(n54), .B(n50), .Z(N100) );
  NR2M1P U44 ( .A(n56), .B(n53), .Z(N111) );
  NR2M1P U45 ( .A(n54), .B(n42), .Z(N112) );
  NR2M1P U46 ( .A(n42), .B(n55), .Z(N113) );
  NR2M1P U47 ( .A(n53), .B(n42), .Z(N115) );
  NR2M1P U48 ( .A(n54), .B(n43), .Z(N116) );
  NR2M1P U49 ( .A(n55), .B(n43), .Z(N117) );
  NR2M1P U50 ( .A(n53), .B(n43), .Z(N119) );
  NR2M1P U51 ( .A(n50), .B(n55), .Z(N101) );
  NR2M1P U52 ( .A(n54), .B(n44), .Z(N120) );
  NR2M1P U53 ( .A(n55), .B(n44), .Z(N121) );
  NR2M1P U54 ( .A(n53), .B(n44), .Z(N123) );
  NR2M1P U55 ( .A(n54), .B(n45), .Z(N124) );
  NR2M1P U56 ( .A(n55), .B(n45), .Z(N125) );
  NR2M1P U57 ( .A(n53), .B(n45), .Z(N127) );
  NR2M1P U58 ( .A(n54), .B(n47), .Z(N128) );
  NR2M1P U59 ( .A(n55), .B(n47), .Z(N129) );
  NR2M1P U60 ( .A(n53), .B(n47), .Z(N131) );
  NR3M1P U61 ( .A(bitCount[4]), .B(n54), .C(n49), .Z(N132) );
  NR2M1P U62 ( .A(n50), .B(n53), .Z(N103) );
  NR2M1P U63 ( .A(n54), .B(n52), .Z(N104) );
  NR2M1P U64 ( .A(n55), .B(n52), .Z(N105) );
  NR2M1P U65 ( .A(n53), .B(n52), .Z(N107) );
  NR2M1P U66 ( .A(n54), .B(n56), .Z(N108) );
  NR2M1P U67 ( .A(n56), .B(n55), .Z(N109) );
  NR2M1P U68 ( .A(bitCount[5]), .B(bitCount[4]), .Z(n51) );
  NR2M1P U69 ( .A(bitCount[2]), .B(bitCount[3]), .Z(n48) );
  ND2M1P U70 ( .A(n51), .B(n48), .Z(n50) );
  ND3M1P U71 ( .A(n51), .B(bitCount[3]), .C(n124), .Z(n56) );
  ND2M1P U72 ( .A(bitCount[1]), .B(bitCount[0]), .Z(n53) );
  ND3M1P U73 ( .A(n51), .B(bitCount[2]), .C(bitCount[3]), .Z(n42) );
  ND3M1P U74 ( .A(bitCount[2]), .B(n46), .C(n57), .Z(n44) );
  ND3M1P U75 ( .A(bitCount[3]), .B(n46), .C(n124), .Z(n45) );
  ND3M1P U76 ( .A(bitCount[2]), .B(bitCount[3]), .C(n46), .Z(n47) );
  ND2M1P U77 ( .A(bitCount[5]), .B(n48), .Z(n49) );
  ND3M1P U78 ( .A(bitCount[2]), .B(n51), .C(n57), .Z(n52) );
  AOI22M1P U79 ( .A(transmissionPacket[5]), .B(N127), .C(transmissionPacket[3]), .D(N129), .Z(n62) );
  AOI22M1P U80 ( .A(transmissionPacket[2]), .B(N130), .C(transmissionPacket[1]), .D(N131), .Z(n61) );
  AOI22M1P U81 ( .A(transmissionPacket[32]), .B(N100), .C(
        transmissionPacket[0]), .D(N132), .Z(n60) );
  AOI22M1P U82 ( .A(transmissionPacket[30]), .B(N102), .C(
        transmissionPacket[31]), .D(N101), .Z(n59) );
  ND4M1P U83 ( .A(n62), .B(n61), .C(n60), .D(n59), .Z(n80) );
  AOI22M1P U84 ( .A(transmissionPacket[29]), .B(N103), .C(
        transmissionPacket[28]), .D(N104), .Z(n66) );
  AOI22M1P U85 ( .A(transmissionPacket[27]), .B(N105), .C(
        transmissionPacket[26]), .D(N106), .Z(n65) );
  AOI22M1P U86 ( .A(transmissionPacket[25]), .B(N107), .C(
        transmissionPacket[24]), .D(N108), .Z(n64) );
  AOI22M1P U87 ( .A(transmissionPacket[23]), .B(N109), .C(
        transmissionPacket[22]), .D(N110), .Z(n63) );
  ND4M1P U88 ( .A(n66), .B(n65), .C(n64), .D(n63), .Z(n79) );
  AOI22M1P U89 ( .A(transmissionPacket[20]), .B(N112), .C(
        transmissionPacket[21]), .D(N111), .Z(n70) );
  AOI22M1P U90 ( .A(transmissionPacket[19]), .B(N113), .C(
        transmissionPacket[18]), .D(N114), .Z(n69) );
  AOI22M1P U91 ( .A(transmissionPacket[17]), .B(N115), .C(
        transmissionPacket[16]), .D(N116), .Z(n68) );
  AOI22M1P U92 ( .A(transmissionPacket[15]), .B(N117), .C(
        transmissionPacket[14]), .D(N118), .Z(n67) );
  AND4M1P U93 ( .A(n70), .B(n69), .C(n68), .D(n67), .Z(n77) );
  AOI22M1P U94 ( .A(transmissionPacket[13]), .B(N119), .C(
        transmissionPacket[12]), .D(N120), .Z(n76) );
  AOI22M1P U95 ( .A(transmissionPacket[11]), .B(N121), .C(
        transmissionPacket[10]), .D(N122), .Z(n75) );
  AOI22M1P U96 ( .A(transmissionPacket[9]), .B(N123), .C(transmissionPacket[8]), .D(N124), .Z(n72) );
  AOI22M1P U97 ( .A(transmissionPacket[4]), .B(N128), .C(transmissionPacket[6]), .D(N126), .Z(n71) );
  ND2M1P U98 ( .A(n72), .B(n71), .Z(n73) );
  AOI21M1P U99 ( .A(N125), .B(transmissionPacket[7]), .C(n73), .Z(n74) );
  ND4M1P U100 ( .A(n77), .B(n76), .C(n75), .D(n74), .Z(n78) );
  NR3M1P U101 ( .A(n80), .B(n79), .C(n78), .Z(n83) );
  N1M1P U102 ( .A(n13), .Z(n138) );
  N1M1P U103 ( .A(bitCount[1]), .Z(n128) );
  N1M1P U104 ( .A(bitCount[4]), .Z(n117) );
  ND4DNM1P U105 ( .D(bitCount[3]), .A(n128), .B(n124), .C(n117), .Z(n85) );
  OAI21M1P U106 ( .A(bitCount[0]), .B(n85), .C(bitCount[5]), .Z(n81) );
  AO21CNM1P U107 ( .A(n138), .B(n81), .C(n5), .Z(n82) );
  OAI211M1P U108 ( .A(n83), .B(n131), .C(n15), .D(n82), .Z(N146) );
  N1M1P U109 ( .A(Tx_Ready), .Z(n135) );
  AO21M1P U110 ( .A(n7), .B(n11), .C(n9), .Z(n84) );
  ND3M1P U111 ( .A(Rx_Ready), .B(n135), .C(n84), .Z(n93) );
  N1M1P U112 ( .A(bitCount[5]), .Z(n116) );
  N1M1P U113 ( .A(bitCount[0]), .Z(n130) );
  OR3M1P U114 ( .A(n85), .B(n116), .C(n130), .Z(n86) );
  AOI21M1P U115 ( .A(n135), .B(n86), .C(TxData_Valid), .Z(n162) );
  N1M1P U116 ( .A(transmissionPacket[0]), .Z(n115) );
  AOI22CDNM1P U117 ( .A(TxData[30]), .B(TxData[31]), .C(TxData[31]), .D(
        TxData[30]), .Z(n106) );
  AOI22CDNM1P U118 ( .A(TxData[24]), .B(TxData[25]), .C(TxData[25]), .D(
        TxData[24]), .Z(n90) );
  AOI22CDNM1P U119 ( .A(TxData[26]), .B(TxData[27]), .C(TxData[27]), .D(
        TxData[26]), .Z(n89) );
  N1M1P U120 ( .A(TxData[28]), .Z(n87) );
  AOI22CDNM1P U121 ( .A(TxData[29]), .B(n87), .C(n87), .D(TxData[29]), .Z(n88)
         );
  EN3M1P U122 ( .A(n90), .B(n89), .C(n88), .Z(n105) );
  AOI22CDNM1P U123 ( .A(TxData[6]), .B(TxData[7]), .C(TxData[7]), .D(TxData[6]), .Z(n103) );
  AOI22CDNM1P U124 ( .A(TxData[0]), .B(TxData[1]), .C(TxData[1]), .D(TxData[0]), .Z(n95) );
  AOI22CDNM1P U125 ( .A(TxData[2]), .B(TxData[3]), .C(TxData[3]), .D(TxData[2]), .Z(n94) );
  N1M1P U126 ( .A(TxData[4]), .Z(n91) );
  AOI22CDNM1P U127 ( .A(TxData[5]), .B(n91), .C(n91), .D(TxData[5]), .Z(n92)
         );
  EN3M1P U128 ( .A(n95), .B(n94), .C(n92), .Z(n102) );
  AOI22CDNM1P U129 ( .A(TxData[15]), .B(TxData[16]), .C(TxData[16]), .D(
        TxData[15]), .Z(n99) );
  AOI22CDNM1P U130 ( .A(TxData[17]), .B(TxData[18]), .C(TxData[18]), .D(
        TxData[17]), .Z(n98) );
  N1M1P U131 ( .A(TxData[19]), .Z(n96) );
  AOI22CDNM1P U132 ( .A(TxData[23]), .B(n96), .C(n96), .D(TxData[23]), .Z(n97)
         );
  EN3M1P U133 ( .A(n99), .B(n98), .C(n97), .Z(n100) );
  EN3M1P U134 ( .A(TxData[22]), .B(TxData[14]), .C(n100), .Z(n101) );
  EN3M1P U135 ( .A(n103), .B(n102), .C(n101), .Z(n104) );
  EN3M1P U136 ( .A(n106), .B(n105), .C(n104), .Z(n113) );
  AOI22CDNM1P U137 ( .A(TxData[12]), .B(TxData[13]), .C(TxData[13]), .D(
        TxData[12]), .Z(n109) );
  AOI22CDNM1P U138 ( .A(TxData[8]), .B(TxData[9]), .C(TxData[9]), .D(TxData[8]), .Z(n108) );
  AOI22CDNM1P U139 ( .A(TxData[10]), .B(TxData[11]), .C(TxData[11]), .D(
        TxData[10]), .Z(n107) );
  EN3M1P U140 ( .A(n109), .B(n108), .C(n107), .Z(n110) );
  EN3M1P U141 ( .A(TxData[20]), .B(TxData[21]), .C(n110), .Z(n112) );
  ND2M1P U142 ( .A(n113), .B(n112), .Z(n111) );
  OAI211M1P U143 ( .A(n113), .B(n112), .C(n111), .D(n16), .Z(n114) );
  OAI21M1P U144 ( .A(n16), .B(n115), .C(n114), .Z(n157) );
  NR2M1P U145 ( .A(bitCount[3]), .B(n131), .Z(n121) );
  NR3M1P U146 ( .A(n130), .B(n128), .C(n124), .Z(n120) );
  OAI21M1P U147 ( .A(n120), .B(n131), .C(n15), .Z(n122) );
  NR2M1P U148 ( .A(n121), .B(n122), .Z(n119) );
  ND3M1P U149 ( .A(bitCount[3]), .B(n133), .C(n120), .Z(n118) );
  OAI22M1P U150 ( .A(n119), .B(n116), .C(n117), .D(n118), .Z(n28) );
  AOI22M1P U151 ( .A(bitCount[4]), .B(n119), .C(n118), .D(n117), .Z(n27) );
  AOI22M1P U152 ( .A(bitCount[3]), .B(n122), .C(n121), .D(n120), .Z(n123) );
  N1M1P U153 ( .A(n123), .Z(n26) );
  N1M1P U154 ( .A(n15), .Z(n139) );
  AOI21M1P U155 ( .A(n130), .B(n133), .C(n139), .Z(n129) );
  OA21M1P U156 ( .A(n131), .B(bitCount[1]), .C(n129), .Z(n126) );
  ND3M1P U157 ( .A(bitCount[0]), .B(bitCount[1]), .C(n133), .Z(n125) );
  AOI22M1P U158 ( .A(bitCount[2]), .B(n126), .C(n125), .D(n124), .Z(n25) );
  ND2M1P U159 ( .A(n133), .B(n128), .Z(n127) );
  OAI22M1P U160 ( .A(n129), .B(n128), .C(n130), .D(n127), .Z(n24) );
  AOI22M1P U161 ( .A(bitCount[0]), .B(n15), .C(n131), .D(n130), .Z(n23) );
  N1M1P U162 ( .A(n2), .Z(n141) );
  ND2M1P U163 ( .A(n142), .B(n141), .Z(n14) );
  NR2M1P U164 ( .A(n139), .B(n5), .Z(n132) );
  AOI211M1P U165 ( .A(n138), .B(n139), .C(n133), .D(n132), .Z(n12) );
  NR2M1P U166 ( .A(n7), .B(n93), .Z(n137) );
  N1M1P U167 ( .A(n11), .Z(n134) );
  OR3M1P U168 ( .A(n11), .B(n7), .C(n93), .Z(n136) );
  OAI211M1P U169 ( .A(n137), .B(n134), .C(n135), .D(n136), .Z(n10) );
  AO21CNM1P U170 ( .A(n9), .B(n136), .C(n135), .Z(n8) );
  AO211M1P U171 ( .A(n7), .B(n93), .C(Tx_Ready), .D(n137), .Z(n6) );
  ND3M1P U172 ( .A(n5), .B(n139), .C(n138), .Z(n140) );
endmodule


module rx_0 ( Clk_s, Rst_n, Core_Rcv_Ready, S_Data, RxData_Valid, RxData, 
        Rx_Ready, Rx_Error );
  output [31:0] RxData;
  input Clk_s, Rst_n, Core_Rcv_Ready, S_Data;
  output RxData_Valid, Rx_Ready, Rx_Error;
  wire   bitStuff, N22, N24, N25, N26, dataRx, bufferFull, N27, N229, N242,
         N243, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n223, n224, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248;
  wire   [2:0] zeroCounter;
  wire   [5:0] receivedCounter;

  FD4QM1P startSeq_reg ( .D(n67), .CP(Clk_s), .SD(Rst_n), .Q(n68) );
  FD4QM1P \receivedPacket_reg[0]  ( .D(n65), .CP(Clk_s), .SD(Rst_n), .Q(n66)
         );
  FD4QM1P \receivedPacket_reg[1]  ( .D(n63), .CP(Clk_s), .SD(Rst_n), .Q(n64)
         );
  FD4QM1P \receivedPacket_reg[2]  ( .D(n61), .CP(Clk_s), .SD(Rst_n), .Q(n62)
         );
  FD4QM1P \receivedPacket_reg[3]  ( .D(n59), .CP(Clk_s), .SD(Rst_n), .Q(n60)
         );
  FD4QM1P \receivedPacket_reg[4]  ( .D(n57), .CP(Clk_s), .SD(Rst_n), .Q(n58)
         );
  FD4QM1P \receivedPacket_reg[5]  ( .D(n55), .CP(Clk_s), .SD(Rst_n), .Q(n56)
         );
  FD4QM1P \receivedPacket_reg[6]  ( .D(n53), .CP(Clk_s), .SD(Rst_n), .Q(n54)
         );
  FD4QM1P \receivedPacket_reg[7]  ( .D(n51), .CP(Clk_s), .SD(Rst_n), .Q(n52)
         );
  FD4QM1P \receivedPacket_reg[8]  ( .D(n49), .CP(Clk_s), .SD(Rst_n), .Q(n50)
         );
  FD4QM1P \receivedPacket_reg[9]  ( .D(n47), .CP(Clk_s), .SD(Rst_n), .Q(n48)
         );
  FD4QM1P \receivedPacket_reg[10]  ( .D(n45), .CP(Clk_s), .SD(Rst_n), .Q(n46)
         );
  FD4QM1P \receivedPacket_reg[11]  ( .D(n43), .CP(Clk_s), .SD(Rst_n), .Q(n44)
         );
  FD4QM1P \receivedPacket_reg[12]  ( .D(n41), .CP(Clk_s), .SD(Rst_n), .Q(n42)
         );
  FD4QM1P \receivedPacket_reg[13]  ( .D(n39), .CP(Clk_s), .SD(Rst_n), .Q(n40)
         );
  FD4QM1P \receivedPacket_reg[14]  ( .D(n37), .CP(Clk_s), .SD(Rst_n), .Q(n38)
         );
  FD4QM1P \receivedPacket_reg[15]  ( .D(n35), .CP(Clk_s), .SD(Rst_n), .Q(n36)
         );
  FD4QM1P \receivedPacket_reg[16]  ( .D(n33), .CP(Clk_s), .SD(Rst_n), .Q(n34)
         );
  FD4QM1P \receivedPacket_reg[17]  ( .D(n31), .CP(Clk_s), .SD(Rst_n), .Q(n32)
         );
  FD4QM1P \receivedPacket_reg[18]  ( .D(n29), .CP(Clk_s), .SD(Rst_n), .Q(n30)
         );
  FD4QM1P \receivedPacket_reg[19]  ( .D(n27), .CP(Clk_s), .SD(Rst_n), .Q(n28)
         );
  FD4QM1P \receivedPacket_reg[20]  ( .D(n25), .CP(Clk_s), .SD(Rst_n), .Q(n26)
         );
  FD4QM1P \receivedPacket_reg[21]  ( .D(n23), .CP(Clk_s), .SD(Rst_n), .Q(n24)
         );
  FD4QM1P \receivedPacket_reg[23]  ( .D(n19), .CP(Clk_s), .SD(Rst_n), .Q(n20)
         );
  FD4QM1P \receivedPacket_reg[24]  ( .D(n17), .CP(Clk_s), .SD(Rst_n), .Q(n18)
         );
  FD4QM1P \receivedPacket_reg[25]  ( .D(n15), .CP(Clk_s), .SD(Rst_n), .Q(n16)
         );
  FD4QM1P \receivedPacket_reg[26]  ( .D(n13), .CP(Clk_s), .SD(Rst_n), .Q(n14)
         );
  FD4QM1P \receivedPacket_reg[29]  ( .D(n7), .CP(Clk_s), .SD(Rst_n), .Q(n8) );
  FD4QM1P \receivedPacket_reg[31]  ( .D(n3), .CP(Clk_s), .SD(Rst_n), .Q(n4) );
  FD4QM1P \receivedPacket_reg[32]  ( .D(n1), .CP(Clk_s), .SD(Rst_n), .Q(n2) );
  FD4QM3P \receivedPacket_reg[22]  ( .D(n21), .CP(Clk_s), .SD(Rst_n), .Q(n22)
         );
  FD4QM3P \receivedPacket_reg[28]  ( .D(n9), .CP(Clk_s), .SD(Rst_n), .Q(n10)
         );
  FD4QM3P \receivedPacket_reg[30]  ( .D(n5), .CP(Clk_s), .SD(Rst_n), .Q(n6) );
  FD4QM3P \receivedPacket_reg[27]  ( .D(n11), .CP(Clk_s), .SD(Rst_n), .Q(n12)
         );
  FD2QM1P \zeroCounter_reg[0]  ( .D(N24), .CP(Clk_s), .CD(Rst_n), .Q(
        zeroCounter[0]) );
  FD2QM1P Rx_Ready_reg ( .D(N27), .CP(Clk_s), .CD(Rst_n), .Q(Rx_Ready) );
  FD2QM1P \zeroCounter_reg[1]  ( .D(N25), .CP(Clk_s), .CD(Rst_n), .Q(
        zeroCounter[1]) );
  FD2QM1P \zeroCounter_reg[2]  ( .D(N26), .CP(Clk_s), .CD(Rst_n), .Q(
        zeroCounter[2]) );
  FD2QM1P bitStuff_reg ( .D(N22), .CP(Clk_s), .CD(Rst_n), .Q(bitStuff) );
  FD2QM1P dataRx_reg ( .D(n224), .CP(Clk_s), .CD(Rst_n), .Q(dataRx) );
  FD2QM1P \receivedCounter_reg[0]  ( .D(n223), .CP(Clk_s), .CD(Rst_n), .Q(
        receivedCounter[0]) );
  FD2QM1P Rx_Error_reg ( .D(N229), .CP(Clk_s), .CD(Rst_n), .Q(Rx_Error) );
  FD2QM1P bufferFull_reg ( .D(N242), .CP(Clk_s), .CD(Rst_n), .Q(bufferFull) );
  FD2QM1P \receivedCounter_reg[1]  ( .D(n73), .CP(Clk_s), .CD(Rst_n), .Q(
        receivedCounter[1]) );
  FD2QM1P \receivedCounter_reg[3]  ( .D(n71), .CP(Clk_s), .CD(Rst_n), .Q(
        receivedCounter[3]) );
  FD2QM1P RxData_Valid_reg ( .D(N243), .CP(Clk_s), .CD(Rst_n), .Q(RxData_Valid) );
  FD2QM1P \receivedCounter_reg[2]  ( .D(n72), .CP(Clk_s), .CD(Rst_n), .Q(
        receivedCounter[2]) );
  FD2QM1P \receivedCounter_reg[4]  ( .D(n70), .CP(Clk_s), .CD(Rst_n), .Q(
        receivedCounter[4]) );
  FD2QM1P \receivedCounter_reg[5]  ( .D(n69), .CP(Clk_s), .CD(Rst_n), .Q(
        receivedCounter[5]) );
  FD2QM1P \RxData_reg[27]  ( .D(n162), .CP(Clk_s), .CD(Rst_n), .Q(RxData[27])
         );
  FD2QM1P \RxData_reg[21]  ( .D(n168), .CP(Clk_s), .CD(Rst_n), .Q(RxData[21])
         );
  FD2QM1P \RxData_reg[22]  ( .D(n167), .CP(Clk_s), .CD(Rst_n), .Q(RxData[22])
         );
  FD2QM1P \RxData_reg[16]  ( .D(n173), .CP(Clk_s), .CD(Rst_n), .Q(RxData[16])
         );
  FD2QM1P \RxData_reg[14]  ( .D(n175), .CP(Clk_s), .CD(Rst_n), .Q(RxData[14])
         );
  FD2QM1P \RxData_reg[10]  ( .D(n179), .CP(Clk_s), .CD(Rst_n), .Q(RxData[10])
         );
  FD2QM1P \RxData_reg[1]  ( .D(n188), .CP(Clk_s), .CD(Rst_n), .Q(RxData[1]) );
  FD2QM1P \RxData_reg[23]  ( .D(n166), .CP(Clk_s), .CD(Rst_n), .Q(RxData[23])
         );
  FD2QM1P \RxData_reg[15]  ( .D(n174), .CP(Clk_s), .CD(Rst_n), .Q(RxData[15])
         );
  FD2QM1P \RxData_reg[6]  ( .D(n183), .CP(Clk_s), .CD(Rst_n), .Q(RxData[6]) );
  FD2QM1P \RxData_reg[5]  ( .D(n184), .CP(Clk_s), .CD(Rst_n), .Q(RxData[5]) );
  FD2QM1P \RxData_reg[29]  ( .D(n160), .CP(Clk_s), .CD(Rst_n), .Q(RxData[29])
         );
  FD2QM1P \RxData_reg[26]  ( .D(n163), .CP(Clk_s), .CD(Rst_n), .Q(RxData[26])
         );
  FD2QM1P \RxData_reg[31]  ( .D(n158), .CP(Clk_s), .CD(Rst_n), .Q(RxData[31])
         );
  FD2QM1P \RxData_reg[24]  ( .D(n165), .CP(Clk_s), .CD(Rst_n), .Q(RxData[24])
         );
  FD2QM1P \RxData_reg[19]  ( .D(n170), .CP(Clk_s), .CD(Rst_n), .Q(RxData[19])
         );
  FD2QM1P \RxData_reg[17]  ( .D(n172), .CP(Clk_s), .CD(Rst_n), .Q(RxData[17])
         );
  FD2QM1P \RxData_reg[13]  ( .D(n176), .CP(Clk_s), .CD(Rst_n), .Q(RxData[13])
         );
  FD2QM1P \RxData_reg[8]  ( .D(n181), .CP(Clk_s), .CD(Rst_n), .Q(RxData[8]) );
  FD2QM1P \RxData_reg[4]  ( .D(n185), .CP(Clk_s), .CD(Rst_n), .Q(RxData[4]) );
  FD2QM1P \RxData_reg[3]  ( .D(n186), .CP(Clk_s), .CD(Rst_n), .Q(RxData[3]) );
  FD2QM1P \RxData_reg[0]  ( .D(n189), .CP(Clk_s), .CD(Rst_n), .Q(RxData[0]) );
  FD2QM1P \RxData_reg[20]  ( .D(n169), .CP(Clk_s), .CD(Rst_n), .Q(RxData[20])
         );
  FD2QM1P \RxData_reg[12]  ( .D(n177), .CP(Clk_s), .CD(Rst_n), .Q(RxData[12])
         );
  FD2QM1P \RxData_reg[9]  ( .D(n180), .CP(Clk_s), .CD(Rst_n), .Q(RxData[9]) );
  FD2QM1P \RxData_reg[2]  ( .D(n187), .CP(Clk_s), .CD(Rst_n), .Q(RxData[2]) );
  FD2QM1P \RxData_reg[30]  ( .D(n159), .CP(Clk_s), .CD(Rst_n), .Q(RxData[30])
         );
  FD2QM1P \RxData_reg[25]  ( .D(n164), .CP(Clk_s), .CD(Rst_n), .Q(RxData[25])
         );
  FD2QM1P \RxData_reg[18]  ( .D(n171), .CP(Clk_s), .CD(Rst_n), .Q(RxData[18])
         );
  FD2QM1P \RxData_reg[11]  ( .D(n178), .CP(Clk_s), .CD(Rst_n), .Q(RxData[11])
         );
  FD2QM1P \RxData_reg[7]  ( .D(n182), .CP(Clk_s), .CD(Rst_n), .Q(RxData[7]) );
  FD2QM1P \RxData_reg[28]  ( .D(n161), .CP(Clk_s), .CD(Rst_n), .Q(RxData[28])
         );
  NR2M2P U3 ( .A(n227), .B(bitStuff), .Z(n119) );
  ND2M1P U4 ( .A(n119), .B(n117), .Z(n77) );
  N1M10P U5 ( .A(n75), .Z(n74) );
  N1M1P U6 ( .A(n12), .Z(n244) );
  N1M1P U7 ( .A(n6), .Z(n247) );
  N1M1P U8 ( .A(n8), .Z(n246) );
  N1M1P U9 ( .A(n10), .Z(n245) );
  N1M2P U10 ( .A(n81), .Z(n80) );
  N1M3P U11 ( .A(n77), .Z(n78) );
  N1M2P U12 ( .A(n81), .Z(n79) );
  AOI22DNM1P U13 ( .A(n154), .B(n78), .D(n2), .C(n79), .Z(n1) );
  N1M6P U14 ( .A(n151), .Z(n75) );
  ND2M1P U15 ( .A(dataRx), .B(n68), .Z(n227) );
  N1M8P U16 ( .A(n75), .Z(n76) );
  ND2FM3P U17 ( .A(n208), .B(n119), .Z(n151) );
  NR2M4P U18 ( .A(n118), .B(n117), .Z(n208) );
  EOFM1P U19 ( .A(n30), .B(n107), .Z(n108) );
  ND2M3P U20 ( .A(n115), .B(n229), .Z(n118) );
  ENM2P U21 ( .A(n114), .B(n113), .Z(n115) );
  OAI21M2P U22 ( .A(n84), .B(n83), .C(receivedCounter[5]), .Z(n117) );
  N1M1P U23 ( .A(bufferFull), .Z(n229) );
  OR2M1P U24 ( .A(receivedCounter[3]), .B(receivedCounter[0]), .Z(n83) );
  NR2BNM1P U25 ( .B(n119), .A(n117), .Z(n116) );
  ND2BNM1P U26 ( .B(receivedCounter[1]), .A(n82), .Z(n84) );
  AOI22M1P U27 ( .A(n154), .B(n80), .C(n247), .D(n78), .Z(n3) );
  N1M1P U28 ( .A(n14), .Z(n215) );
  N1M1P U29 ( .A(n16), .Z(n214) );
  N1M1P U30 ( .A(n20), .Z(n212) );
  N1M1P U31 ( .A(n22), .Z(n211) );
  AOI22M1P U32 ( .A(n210), .B(n80), .C(n78), .D(n155), .Z(n23) );
  N1M1P U33 ( .A(n24), .Z(n210) );
  OAI21M1P U34 ( .A(n229), .B(n222), .C(n209), .Z(N242) );
  N1M1P U35 ( .A(receivedCounter[3]), .Z(n218) );
  AOI22M1P U36 ( .A(n207), .B(n79), .C(n243), .D(S_Data), .Z(n65) );
  N1M1P U37 ( .A(receivedCounter[4]), .Z(n217) );
  N1M1P U38 ( .A(receivedCounter[0]), .Z(n216) );
  N1M1P U39 ( .A(receivedCounter[2]), .Z(n219) );
  AOI22M1P U40 ( .A(n204), .B(n79), .C(n78), .D(n205), .Z(n59) );
  AOI22M1P U41 ( .A(n195), .B(n79), .C(n78), .D(n196), .Z(n41) );
  AOI22M1P U42 ( .A(n193), .B(n79), .C(n78), .D(n194), .Z(n37) );
  AOI22M1P U43 ( .A(n197), .B(n79), .C(n78), .D(n198), .Z(n45) );
  AOI22M1P U44 ( .A(n199), .B(n79), .C(n78), .D(n200), .Z(n49) );
  AOI22M1P U45 ( .A(n196), .B(n79), .C(n78), .D(n197), .Z(n43) );
  N1M1P U46 ( .A(n46), .Z(n197) );
  N1M1P U47 ( .A(n44), .Z(n196) );
  AOI22M1P U48 ( .A(n200), .B(n79), .C(n78), .D(n201), .Z(n51) );
  N1M1P U49 ( .A(n52), .Z(n200) );
  AOI22M1P U50 ( .A(n201), .B(n79), .C(n78), .D(n202), .Z(n53) );
  N1M1P U51 ( .A(n54), .Z(n201) );
  AOI22M1P U52 ( .A(n190), .B(n79), .C(n78), .D(n191), .Z(n31) );
  AOI22M1P U53 ( .A(n202), .B(n79), .C(n78), .D(n203), .Z(n55) );
  N1M1P U54 ( .A(n56), .Z(n202) );
  AOI22M1P U55 ( .A(n203), .B(n79), .C(n78), .D(n204), .Z(n57) );
  N1M1P U56 ( .A(n60), .Z(n204) );
  N1M1P U57 ( .A(n58), .Z(n203) );
  AOI22M1P U58 ( .A(n194), .B(n79), .C(n78), .D(n195), .Z(n39) );
  N1M1P U59 ( .A(n42), .Z(n195) );
  N1M1P U60 ( .A(n40), .Z(n194) );
  AOI22M1P U61 ( .A(n205), .B(n79), .C(n78), .D(n206), .Z(n61) );
  N1M1P U62 ( .A(n62), .Z(n205) );
  N1M1P U63 ( .A(n4), .Z(n154) );
  AOI22M1P U64 ( .A(n157), .B(n79), .C(n78), .D(n190), .Z(n29) );
  N1M1P U65 ( .A(n32), .Z(n190) );
  AOI22M1P U66 ( .A(n155), .B(n79), .C(n78), .D(n156), .Z(n25) );
  N1M1P U67 ( .A(n26), .Z(n155) );
  AOI22M1P U68 ( .A(n191), .B(n79), .C(n78), .D(n192), .Z(n33) );
  N1M1P U69 ( .A(n34), .Z(n191) );
  AOI22M1P U70 ( .A(n156), .B(n79), .C(n78), .D(n157), .Z(n27) );
  N1M1P U71 ( .A(n28), .Z(n156) );
  AOI22M1P U72 ( .A(n192), .B(n79), .C(n78), .D(n193), .Z(n35) );
  N1M1P U73 ( .A(n38), .Z(n193) );
  N1M1P U74 ( .A(n36), .Z(n192) );
  AOI22M1P U75 ( .A(n198), .B(n79), .C(n78), .D(n199), .Z(n47) );
  N1M1P U76 ( .A(n50), .Z(n199) );
  N1M1P U77 ( .A(n48), .Z(n198) );
  AOI22M1P U78 ( .A(n206), .B(n79), .C(n78), .D(n207), .Z(n63) );
  N1M1P U79 ( .A(n66), .Z(n207) );
  ND2BNM1P U80 ( .B(n229), .A(n116), .Z(n85) );
  N1M1P U81 ( .A(n64), .Z(n206) );
  MUX21LM1P U82 ( .A(n18), .B(n143), .S(n76), .Z(n166) );
  N1M1P U83 ( .A(RxData[23]), .Z(n143) );
  MUX21LM1P U84 ( .A(n10), .B(n147), .S(n76), .Z(n162) );
  N1M1P U85 ( .A(RxData[27]), .Z(n147) );
  MUX21LM1P U86 ( .A(n12), .B(n146), .S(n74), .Z(n163) );
  N1M1P U87 ( .A(RxData[26]), .Z(n146) );
  MUX21LM1P U88 ( .A(n8), .B(n148), .S(n74), .Z(n161) );
  N1M1P U89 ( .A(RxData[28]), .Z(n148) );
  MUX21LM1P U90 ( .A(n16), .B(n144), .S(n74), .Z(n165) );
  N1M1P U91 ( .A(RxData[24]), .Z(n144) );
  MUX21LM1P U92 ( .A(n2), .B(n152), .S(n74), .Z(n158) );
  N1M1P U93 ( .A(RxData[31]), .Z(n152) );
  MUX21LM1P U94 ( .A(n20), .B(n142), .S(n76), .Z(n167) );
  N1M1P U95 ( .A(RxData[22]), .Z(n142) );
  MUX21LM1P U96 ( .A(n6), .B(n149), .S(n74), .Z(n160) );
  N1M1P U97 ( .A(RxData[29]), .Z(n149) );
  MUX21LM1P U98 ( .A(n14), .B(n145), .S(n74), .Z(n164) );
  N1M1P U99 ( .A(RxData[25]), .Z(n145) );
  MUX21LM1P U100 ( .A(n4), .B(n150), .S(n74), .Z(n159) );
  N1M1P U101 ( .A(RxData[30]), .Z(n150) );
  MUX21LM1P U102 ( .A(n30), .B(n137), .S(n74), .Z(n172) );
  N1M1P U103 ( .A(RxData[17]), .Z(n137) );
  MUX21LM1P U104 ( .A(n22), .B(n141), .S(n76), .Z(n168) );
  N1M1P U105 ( .A(RxData[21]), .Z(n141) );
  MUX21LM1P U106 ( .A(n62), .B(n121), .S(n76), .Z(n188) );
  N1M1P U107 ( .A(RxData[1]), .Z(n121) );
  MUX21LM1P U108 ( .A(n26), .B(n139), .S(n74), .Z(n170) );
  N1M1P U109 ( .A(RxData[19]), .Z(n139) );
  MUX21LM1P U110 ( .A(n36), .B(n134), .S(n76), .Z(n175) );
  N1M1P U111 ( .A(RxData[14]), .Z(n134) );
  MUX21LM1P U112 ( .A(n32), .B(n136), .S(n76), .Z(n173) );
  N1M1P U113 ( .A(RxData[16]), .Z(n136) );
  MUX21LM1P U114 ( .A(n48), .B(n128), .S(n74), .Z(n181) );
  N1M1P U115 ( .A(RxData[8]), .Z(n128) );
  MUX21LM1P U116 ( .A(n56), .B(n124), .S(n74), .Z(n185) );
  N1M1P U117 ( .A(RxData[4]), .Z(n124) );
  MUX21LM1P U118 ( .A(n38), .B(n133), .S(n74), .Z(n176) );
  N1M1P U119 ( .A(RxData[13]), .Z(n133) );
  MUX21LM1P U120 ( .A(n64), .B(n120), .S(n74), .Z(n189) );
  N1M1P U121 ( .A(RxData[0]), .Z(n120) );
  MUX21LM1P U122 ( .A(n58), .B(n123), .S(n74), .Z(n186) );
  N1M1P U123 ( .A(RxData[3]), .Z(n123) );
  MUX21LM1P U124 ( .A(n44), .B(n130), .S(n76), .Z(n179) );
  N1M1P U125 ( .A(RxData[10]), .Z(n130) );
  MUX21LM1P U126 ( .A(n46), .B(n129), .S(n74), .Z(n180) );
  N1M1P U127 ( .A(RxData[9]), .Z(n129) );
  MUX21LM1P U128 ( .A(n24), .B(n140), .S(n74), .Z(n169) );
  N1M1P U129 ( .A(RxData[20]), .Z(n140) );
  MUX21LM1P U130 ( .A(n60), .B(n122), .S(n74), .Z(n187) );
  N1M1P U131 ( .A(RxData[2]), .Z(n122) );
  MUX21LM1P U132 ( .A(n34), .B(n135), .S(n76), .Z(n174) );
  N1M1P U133 ( .A(RxData[15]), .Z(n135) );
  MUX21LM1P U134 ( .A(n40), .B(n132), .S(n74), .Z(n177) );
  N1M1P U135 ( .A(RxData[12]), .Z(n132) );
  MUX21LM1P U136 ( .A(n54), .B(n125), .S(n76), .Z(n184) );
  N1M1P U137 ( .A(RxData[5]), .Z(n125) );
  MUX21LM1P U138 ( .A(n52), .B(n126), .S(n76), .Z(n183) );
  N1M1P U139 ( .A(RxData[6]), .Z(n126) );
  MUX21LM1P U140 ( .A(n42), .B(n131), .S(n74), .Z(n178) );
  N1M1P U141 ( .A(RxData[11]), .Z(n131) );
  MUX21LM1P U142 ( .A(n50), .B(n127), .S(n74), .Z(n182) );
  N1M1P U143 ( .A(RxData[7]), .Z(n127) );
  MUX21LM1P U144 ( .A(n28), .B(n138), .S(n74), .Z(n171) );
  NR2M1P U145 ( .A(receivedCounter[2]), .B(receivedCounter[4]), .Z(n82) );
  ENFM1P U146 ( .A(n112), .B(n111), .Z(n113) );
  EOFM1P U147 ( .A(n110), .B(n109), .Z(n111) );
  EOFM1P U148 ( .A(n221), .B(n108), .Z(n109) );
  N1M1P U149 ( .A(n30), .Z(n157) );
  AOI22M1P U150 ( .A(n6), .B(n8), .C(n246), .D(n247), .Z(n221) );
  EOFM1P U151 ( .A(n26), .B(n28), .Z(n106) );
  ENFM1P U152 ( .A(n105), .B(n104), .Z(n112) );
  ENFM1P U153 ( .A(n103), .B(n102), .Z(n104) );
  ENFM1P U154 ( .A(n32), .B(n34), .Z(n102) );
  ENFM1P U155 ( .A(n36), .B(n54), .Z(n103) );
  ENFM1P U156 ( .A(n101), .B(n100), .Z(n105) );
  EOFM1P U157 ( .A(n56), .B(n42), .Z(n100) );
  ENFM1P U158 ( .A(n44), .B(n46), .Z(n101) );
  ENFM1P U159 ( .A(n99), .B(n98), .Z(n114) );
  ENFM1P U160 ( .A(n97), .B(n96), .Z(n98) );
  ENFM1P U161 ( .A(n95), .B(n94), .Z(n96) );
  EOFM1P U162 ( .A(n48), .B(n50), .Z(n94) );
  ENFM1P U163 ( .A(n58), .B(n52), .Z(n95) );
  ENFM1P U164 ( .A(n93), .B(n92), .Z(n97) );
  EOFM1P U165 ( .A(n62), .B(n4), .Z(n92) );
  ENFM1P U166 ( .A(n64), .B(n60), .Z(n93) );
  ENFM1P U167 ( .A(n91), .B(n90), .Z(n99) );
  ENFM1P U168 ( .A(n89), .B(n88), .Z(n90) );
  ENFM1P U169 ( .A(n38), .B(n40), .Z(n88) );
  ENFM1P U170 ( .A(n2), .B(n66), .Z(n89) );
  ENFM1P U171 ( .A(n87), .B(n86), .Z(n91) );
  ENFM1P U172 ( .A(n16), .B(n24), .Z(n86) );
  EOFM1P U173 ( .A(n20), .B(n14), .Z(n87) );
  N1M1P U174 ( .A(RxData[18]), .Z(n138) );
  N1M2P U175 ( .A(n248), .Z(n81) );
  OAI21M1P U176 ( .A(n227), .B(n228), .C(n85), .Z(n248) );
  N1M1P U177 ( .A(n18), .Z(n213) );
  AND3M1P U178 ( .A(n118), .B(n116), .C(n229), .Z(N229) );
  ENFM1P U179 ( .A(n22), .B(n18), .Z(n107) );
  N1M1P U180 ( .A(n208), .Z(n209) );
  NR2BNM1P U181 ( .B(RxData_Valid), .A(n208), .Z(n153) );
  EOFM1P U182 ( .A(n106), .B(n220), .Z(n110) );
  OA21M1P U183 ( .A(n153), .B(bufferFull), .C(Core_Rcv_Ready), .Z(N243) );
  ND2M1P U184 ( .A(zeroCounter[1]), .B(zeroCounter[0]), .Z(n225) );
  NR3M1P U185 ( .A(S_Data), .B(zeroCounter[2]), .C(n225), .Z(N26) );
  N1M1P U186 ( .A(receivedCounter[5]), .Z(n241) );
  AND2M1P U187 ( .A(N26), .B(n241), .Z(N22) );
  AOI22M1P U188 ( .A(n10), .B(n12), .C(n244), .D(n245), .Z(n220) );
  NR3M1P U189 ( .A(S_Data), .B(zeroCounter[2]), .C(zeroCounter[0]), .Z(N24) );
  NR2BNM1P U190 ( .B(RxData_Valid), .A(Core_Rcv_Ready), .Z(n222) );
  OAI21M1P U191 ( .A(zeroCounter[1]), .B(zeroCounter[0]), .C(n225), .Z(n226)
         );
  NR3M1P U192 ( .A(S_Data), .B(zeroCounter[2]), .C(n226), .Z(N25) );
  NR2BNM1P U193 ( .B(n68), .A(dataRx), .Z(N27) );
  ND2M1P U194 ( .A(n68), .B(n77), .Z(n243) );
  N1M1P U195 ( .A(bitStuff), .Z(n228) );
  ND2BNM1P U196 ( .B(n243), .A(n81), .Z(n224) );
  ND2M1P U197 ( .A(n78), .B(n216), .Z(n230) );
  OAI211M1P U198 ( .A(n81), .B(n216), .C(n68), .D(n230), .Z(n223) );
  AOI21M1P U199 ( .A(n78), .B(n216), .C(n80), .Z(n231) );
  N1M1P U200 ( .A(receivedCounter[1]), .Z(n235) );
  NR2M1P U201 ( .A(receivedCounter[1]), .B(n77), .Z(n232) );
  OAI22CDNM1P U202 ( .A(n231), .B(n235), .C(receivedCounter[0]), .D(n232), .Z(
        n73) );
  AOI211M1P U203 ( .A(n78), .B(n216), .C(n232), .D(n80), .Z(n234) );
  ND3M1P U204 ( .A(receivedCounter[1]), .B(receivedCounter[0]), .C(n78), .Z(
        n233) );
  AOI22M1P U205 ( .A(receivedCounter[2]), .B(n234), .C(n233), .D(n219), .Z(n72) );
  NR3M1P U206 ( .A(n235), .B(n219), .C(n216), .Z(n239) );
  N1M1P U207 ( .A(n239), .Z(n236) );
  AOI21M1P U208 ( .A(n236), .B(n78), .C(n80), .Z(n238) );
  ND2M1P U209 ( .A(n78), .B(n218), .Z(n237) );
  OAI22M1P U210 ( .A(n238), .B(n218), .C(n237), .D(n236), .Z(n71) );
  OA21M1P U211 ( .A(n77), .B(receivedCounter[3]), .C(n238), .Z(n242) );
  ND3M1P U212 ( .A(receivedCounter[3]), .B(n78), .C(n239), .Z(n240) );
  AOI22M1P U213 ( .A(receivedCounter[4]), .B(n242), .C(n240), .D(n217), .Z(n70) );
  OAI22M1P U214 ( .A(n242), .B(n241), .C(n217), .D(n240), .Z(n69) );
  ND2BNM1P U215 ( .B(S_Data), .A(zeroCounter[2]), .Z(n67) );
  AOI22M1P U216 ( .A(n78), .B(n210), .C(n211), .D(n80), .Z(n21) );
  AOI22M1P U217 ( .A(n78), .B(n211), .C(n212), .D(n80), .Z(n19) );
  AOI22M1P U218 ( .A(n78), .B(n212), .C(n213), .D(n80), .Z(n17) );
  AOI22M1P U219 ( .A(n78), .B(n213), .C(n214), .D(n80), .Z(n15) );
  AOI22M1P U220 ( .A(n78), .B(n214), .C(n215), .D(n80), .Z(n13) );
  AOI22M1P U221 ( .A(n78), .B(n215), .C(n244), .D(n80), .Z(n11) );
  AOI22M1P U222 ( .A(n78), .B(n244), .C(n245), .D(n80), .Z(n9) );
  AOI22M1P U223 ( .A(n78), .B(n245), .C(n246), .D(n80), .Z(n7) );
  AOI22M1P U224 ( .A(n78), .B(n246), .C(n247), .D(n80), .Z(n5) );
endmodule


module rx_1 ( Clk_s, Rst_n, Core_Rcv_Ready, S_Data, RxData_Valid, RxData, 
        Rx_Ready, Rx_Error );
  output [31:0] RxData;
  input Clk_s, Rst_n, Core_Rcv_Ready, S_Data;
  output RxData_Valid, Rx_Ready, Rx_Error;
  wire   bitStuff, N22, N24, N25, N26, dataRx, bufferFull, N27, N229, N242,
         N243, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354;
  wire   [2:0] zeroCounter;
  wire   [5:0] receivedCounter;

  FD4QM1P startSeq_reg ( .D(n288), .CP(Clk_s), .SD(Rst_n), .Q(n287) );
  FD4QM1P \receivedPacket_reg[0]  ( .D(n290), .CP(Clk_s), .SD(Rst_n), .Q(n289)
         );
  FD4QM1P \receivedPacket_reg[1]  ( .D(n292), .CP(Clk_s), .SD(Rst_n), .Q(n291)
         );
  FD4QM1P \receivedPacket_reg[2]  ( .D(n294), .CP(Clk_s), .SD(Rst_n), .Q(n293)
         );
  FD4QM1P \receivedPacket_reg[3]  ( .D(n296), .CP(Clk_s), .SD(Rst_n), .Q(n295)
         );
  FD4QM1P \receivedPacket_reg[4]  ( .D(n298), .CP(Clk_s), .SD(Rst_n), .Q(n297)
         );
  FD4QM1P \receivedPacket_reg[5]  ( .D(n300), .CP(Clk_s), .SD(Rst_n), .Q(n299)
         );
  FD4QM1P \receivedPacket_reg[6]  ( .D(n302), .CP(Clk_s), .SD(Rst_n), .Q(n301)
         );
  FD4QM1P \receivedPacket_reg[7]  ( .D(n304), .CP(Clk_s), .SD(Rst_n), .Q(n303)
         );
  FD4QM1P \receivedPacket_reg[8]  ( .D(n306), .CP(Clk_s), .SD(Rst_n), .Q(n305)
         );
  FD4QM1P \receivedPacket_reg[9]  ( .D(n308), .CP(Clk_s), .SD(Rst_n), .Q(n307)
         );
  FD4QM1P \receivedPacket_reg[10]  ( .D(n310), .CP(Clk_s), .SD(Rst_n), .Q(n309) );
  FD4QM1P \receivedPacket_reg[11]  ( .D(n312), .CP(Clk_s), .SD(Rst_n), .Q(n311) );
  FD4QM1P \receivedPacket_reg[12]  ( .D(n314), .CP(Clk_s), .SD(Rst_n), .Q(n313) );
  FD4QM1P \receivedPacket_reg[13]  ( .D(n316), .CP(Clk_s), .SD(Rst_n), .Q(n315) );
  FD4QM1P \receivedPacket_reg[14]  ( .D(n318), .CP(Clk_s), .SD(Rst_n), .Q(n317) );
  FD4QM1P \receivedPacket_reg[15]  ( .D(n320), .CP(Clk_s), .SD(Rst_n), .Q(n319) );
  FD4QM1P \receivedPacket_reg[16]  ( .D(n322), .CP(Clk_s), .SD(Rst_n), .Q(n321) );
  FD4QM1P \receivedPacket_reg[17]  ( .D(n324), .CP(Clk_s), .SD(Rst_n), .Q(n323) );
  FD4QM1P \receivedPacket_reg[18]  ( .D(n326), .CP(Clk_s), .SD(Rst_n), .Q(n325) );
  FD4QM1P \receivedPacket_reg[19]  ( .D(n328), .CP(Clk_s), .SD(Rst_n), .Q(n327) );
  FD4QM1P \receivedPacket_reg[20]  ( .D(n330), .CP(Clk_s), .SD(Rst_n), .Q(n329) );
  FD4QM1P \receivedPacket_reg[21]  ( .D(n332), .CP(Clk_s), .SD(Rst_n), .Q(n331) );
  FD4QM1P \receivedPacket_reg[24]  ( .D(n338), .CP(Clk_s), .SD(Rst_n), .Q(n337) );
  FD4QM1P \receivedPacket_reg[25]  ( .D(n340), .CP(Clk_s), .SD(Rst_n), .Q(n339) );
  FD4QM1P \receivedPacket_reg[26]  ( .D(n342), .CP(Clk_s), .SD(Rst_n), .Q(n341) );
  FD4QM1P \receivedPacket_reg[29]  ( .D(n348), .CP(Clk_s), .SD(Rst_n), .Q(n347) );
  FD4QM1P \receivedPacket_reg[31]  ( .D(n352), .CP(Clk_s), .SD(Rst_n), .Q(n351) );
  FD4QM1P \receivedPacket_reg[32]  ( .D(n354), .CP(Clk_s), .SD(Rst_n), .Q(n353) );
  FD2QM1P \RxData_reg[31]  ( .D(n281), .CP(Clk_s), .CD(Rst_n), .Q(RxData[31])
         );
  FD2QM1P \RxData_reg[30]  ( .D(n280), .CP(Clk_s), .CD(Rst_n), .Q(RxData[30])
         );
  FD2QM1P \RxData_reg[29]  ( .D(n279), .CP(Clk_s), .CD(Rst_n), .Q(RxData[29])
         );
  FD2QM1P \RxData_reg[28]  ( .D(n278), .CP(Clk_s), .CD(Rst_n), .Q(RxData[28])
         );
  FD2QM1P \RxData_reg[27]  ( .D(n277), .CP(Clk_s), .CD(Rst_n), .Q(RxData[27])
         );
  FD2QM1P \RxData_reg[26]  ( .D(n276), .CP(Clk_s), .CD(Rst_n), .Q(RxData[26])
         );
  FD2QM1P \RxData_reg[25]  ( .D(n275), .CP(Clk_s), .CD(Rst_n), .Q(RxData[25])
         );
  FD2QM1P \RxData_reg[24]  ( .D(n274), .CP(Clk_s), .CD(Rst_n), .Q(RxData[24])
         );
  FD2QM1P \RxData_reg[23]  ( .D(n273), .CP(Clk_s), .CD(Rst_n), .Q(RxData[23])
         );
  FD2QM1P \RxData_reg[22]  ( .D(n272), .CP(Clk_s), .CD(Rst_n), .Q(RxData[22])
         );
  FD2QM1P \RxData_reg[21]  ( .D(n271), .CP(Clk_s), .CD(Rst_n), .Q(RxData[21])
         );
  FD2QM1P \RxData_reg[20]  ( .D(n270), .CP(Clk_s), .CD(Rst_n), .Q(RxData[20])
         );
  FD2QM1P \RxData_reg[19]  ( .D(n269), .CP(Clk_s), .CD(Rst_n), .Q(RxData[19])
         );
  FD2QM1P \RxData_reg[18]  ( .D(n268), .CP(Clk_s), .CD(Rst_n), .Q(RxData[18])
         );
  FD2QM1P \RxData_reg[17]  ( .D(n267), .CP(Clk_s), .CD(Rst_n), .Q(RxData[17])
         );
  FD2QM1P \RxData_reg[16]  ( .D(n266), .CP(Clk_s), .CD(Rst_n), .Q(RxData[16])
         );
  FD2QM1P \RxData_reg[15]  ( .D(n265), .CP(Clk_s), .CD(Rst_n), .Q(RxData[15])
         );
  FD2QM1P \RxData_reg[14]  ( .D(n264), .CP(Clk_s), .CD(Rst_n), .Q(RxData[14])
         );
  FD2QM1P \RxData_reg[13]  ( .D(n263), .CP(Clk_s), .CD(Rst_n), .Q(RxData[13])
         );
  FD2QM1P \RxData_reg[12]  ( .D(n262), .CP(Clk_s), .CD(Rst_n), .Q(RxData[12])
         );
  FD2QM1P \RxData_reg[11]  ( .D(n261), .CP(Clk_s), .CD(Rst_n), .Q(RxData[11])
         );
  FD2QM1P \RxData_reg[10]  ( .D(n260), .CP(Clk_s), .CD(Rst_n), .Q(RxData[10])
         );
  FD2QM1P \RxData_reg[9]  ( .D(n259), .CP(Clk_s), .CD(Rst_n), .Q(RxData[9]) );
  FD2QM1P \RxData_reg[8]  ( .D(n258), .CP(Clk_s), .CD(Rst_n), .Q(RxData[8]) );
  FD2QM1P \RxData_reg[7]  ( .D(n257), .CP(Clk_s), .CD(Rst_n), .Q(RxData[7]) );
  FD2QM1P \RxData_reg[6]  ( .D(n256), .CP(Clk_s), .CD(Rst_n), .Q(RxData[6]) );
  FD2QM1P \RxData_reg[5]  ( .D(n255), .CP(Clk_s), .CD(Rst_n), .Q(RxData[5]) );
  FD2QM1P \RxData_reg[4]  ( .D(n254), .CP(Clk_s), .CD(Rst_n), .Q(RxData[4]) );
  FD2QM1P \RxData_reg[3]  ( .D(n253), .CP(Clk_s), .CD(Rst_n), .Q(RxData[3]) );
  FD2QM1P \RxData_reg[2]  ( .D(n252), .CP(Clk_s), .CD(Rst_n), .Q(RxData[2]) );
  FD2QM1P \RxData_reg[1]  ( .D(n251), .CP(Clk_s), .CD(Rst_n), .Q(RxData[1]) );
  FD2QM1P \RxData_reg[0]  ( .D(n250), .CP(Clk_s), .CD(Rst_n), .Q(RxData[0]) );
  FD4QM3P \receivedPacket_reg[28]  ( .D(n346), .CP(Clk_s), .SD(Rst_n), .Q(n345) );
  FD4QM3P \receivedPacket_reg[27]  ( .D(n344), .CP(Clk_s), .SD(Rst_n), .Q(n343) );
  FD4QM3P \receivedPacket_reg[22]  ( .D(n334), .CP(Clk_s), .SD(Rst_n), .Q(n333) );
  FD2QM1P \zeroCounter_reg[0]  ( .D(N24), .CP(Clk_s), .CD(Rst_n), .Q(
        zeroCounter[0]) );
  FD2QM1P Rx_Ready_reg ( .D(N27), .CP(Clk_s), .CD(Rst_n), .Q(Rx_Ready) );
  FD2QM1P \zeroCounter_reg[1]  ( .D(N25), .CP(Clk_s), .CD(Rst_n), .Q(
        zeroCounter[1]) );
  FD2QM1P \zeroCounter_reg[2]  ( .D(N26), .CP(Clk_s), .CD(Rst_n), .Q(
        zeroCounter[2]) );
  FD2QM1P bitStuff_reg ( .D(N22), .CP(Clk_s), .CD(Rst_n), .Q(bitStuff) );
  FD2QM1P dataRx_reg ( .D(n248), .CP(Clk_s), .CD(Rst_n), .Q(dataRx) );
  FD2QM1P \receivedCounter_reg[0]  ( .D(n249), .CP(Clk_s), .CD(Rst_n), .Q(
        receivedCounter[0]) );
  FD2QM1P Rx_Error_reg ( .D(N229), .CP(Clk_s), .CD(Rst_n), .Q(Rx_Error) );
  FD2QM1P bufferFull_reg ( .D(N242), .CP(Clk_s), .CD(Rst_n), .Q(bufferFull) );
  FD2QM1P \receivedCounter_reg[1]  ( .D(n282), .CP(Clk_s), .CD(Rst_n), .Q(
        receivedCounter[1]) );
  FD2QM1P \receivedCounter_reg[3]  ( .D(n284), .CP(Clk_s), .CD(Rst_n), .Q(
        receivedCounter[3]) );
  FD2QM1P RxData_Valid_reg ( .D(N243), .CP(Clk_s), .CD(Rst_n), .Q(RxData_Valid) );
  FD2QM1P \receivedCounter_reg[2]  ( .D(n283), .CP(Clk_s), .CD(Rst_n), .Q(
        receivedCounter[2]) );
  FD2QM1P \receivedCounter_reg[4]  ( .D(n285), .CP(Clk_s), .CD(Rst_n), .Q(
        receivedCounter[4]) );
  FD2QM1P \receivedCounter_reg[5]  ( .D(n286), .CP(Clk_s), .CD(Rst_n), .Q(
        receivedCounter[5]) );
  FD4QM1P \receivedPacket_reg[30]  ( .D(n350), .CP(Clk_s), .SD(Rst_n), .Q(n349) );
  FD4QM1P \receivedPacket_reg[23]  ( .D(n336), .CP(Clk_s), .SD(Rst_n), .Q(n335) );
  NR2M2P U3 ( .A(n226), .B(bitStuff), .Z(n118) );
  ND2M1P U4 ( .A(n118), .B(n116), .Z(n78) );
  N1M10P U5 ( .A(n76), .Z(n75) );
  N1M1P U6 ( .A(n347), .Z(n245) );
  N1M1P U7 ( .A(n345), .Z(n244) );
  N1M2P U8 ( .A(n82), .Z(n81) );
  N1M3P U9 ( .A(n78), .Z(n79) );
  N1M2P U10 ( .A(n82), .Z(n80) );
  ENFM1P U11 ( .A(n311), .B(n309), .Z(n74) );
  EN3M1P U12 ( .A(n313), .B(n299), .C(n74), .Z(n104) );
  AOI22DNM1P U13 ( .A(n153), .B(n79), .D(n353), .C(n80), .Z(n354) );
  ND2M3P U14 ( .A(n114), .B(n228), .Z(n117) );
  ND2M1P U15 ( .A(dataRx), .B(n287), .Z(n226) );
  N1M6P U16 ( .A(n150), .Z(n76) );
  N1M6P U17 ( .A(n76), .Z(n77) );
  ND2FM3P U18 ( .A(n207), .B(n118), .Z(n150) );
  ENM2P U19 ( .A(n113), .B(n112), .Z(n114) );
  NR2M4P U20 ( .A(n117), .B(n116), .Z(n207) );
  N1M2P U21 ( .A(n349), .Z(n246) );
  OAI21M2P U22 ( .A(n85), .B(n84), .C(receivedCounter[5]), .Z(n116) );
  N1M1P U23 ( .A(n343), .Z(n243) );
  N1M1P U24 ( .A(bufferFull), .Z(n228) );
  OR2M1P U25 ( .A(receivedCounter[3]), .B(receivedCounter[0]), .Z(n84) );
  NR2BNM1P U26 ( .B(n118), .A(n116), .Z(n115) );
  ND2BNM1P U27 ( .B(receivedCounter[1]), .A(n83), .Z(n85) );
  AND3M1P U28 ( .A(n117), .B(n115), .C(n228), .Z(N229) );
  AOI22M1P U29 ( .A(n153), .B(n81), .C(n246), .D(n79), .Z(n352) );
  N1M1P U30 ( .A(n333), .Z(n210) );
  N1M1P U31 ( .A(n335), .Z(n211) );
  N1M1P U32 ( .A(n337), .Z(n212) );
  N1M1P U33 ( .A(n341), .Z(n214) );
  N1M1P U34 ( .A(n339), .Z(n213) );
  AOI22M1P U35 ( .A(n209), .B(n81), .C(n79), .D(n154), .Z(n332) );
  N1M1P U36 ( .A(n331), .Z(n209) );
  OAI21M1P U37 ( .A(n228), .B(n221), .C(n208), .Z(N242) );
  N1M1P U38 ( .A(n207), .Z(n208) );
  NR2BNM1P U39 ( .B(RxData_Valid), .A(n207), .Z(n152) );
  N1M1P U40 ( .A(receivedCounter[3]), .Z(n217) );
  AOI22M1P U41 ( .A(n206), .B(n80), .C(n242), .D(S_Data), .Z(n290) );
  AOI22M1P U42 ( .A(n199), .B(n80), .C(n79), .D(n200), .Z(n304) );
  AOI22M1P U43 ( .A(n195), .B(n80), .C(n79), .D(n196), .Z(n312) );
  AOI22M1P U44 ( .A(n200), .B(n80), .C(n79), .D(n201), .Z(n302) );
  N1M1P U45 ( .A(n301), .Z(n200) );
  AOI22M1P U46 ( .A(n197), .B(n80), .C(n79), .D(n198), .Z(n308) );
  AOI22M1P U47 ( .A(n201), .B(n80), .C(n79), .D(n202), .Z(n300) );
  N1M1P U48 ( .A(n299), .Z(n201) );
  AOI22M1P U49 ( .A(n191), .B(n80), .C(n79), .D(n192), .Z(n320) );
  AOI22M1P U50 ( .A(n196), .B(n80), .C(n79), .D(n197), .Z(n310) );
  N1M1P U51 ( .A(n307), .Z(n197) );
  N1M1P U52 ( .A(n309), .Z(n196) );
  AOI22M1P U53 ( .A(n202), .B(n80), .C(n79), .D(n203), .Z(n298) );
  N1M1P U54 ( .A(n297), .Z(n202) );
  AOI22M1P U55 ( .A(n155), .B(n80), .C(n79), .D(n156), .Z(n328) );
  AOI22M1P U56 ( .A(n193), .B(n80), .C(n79), .D(n194), .Z(n316) );
  AOI22M1P U57 ( .A(n203), .B(n80), .C(n79), .D(n204), .Z(n296) );
  N1M1P U58 ( .A(n295), .Z(n203) );
  AOI22M1P U59 ( .A(n194), .B(n80), .C(n79), .D(n195), .Z(n314) );
  N1M1P U60 ( .A(n311), .Z(n195) );
  N1M1P U61 ( .A(n313), .Z(n194) );
  AOI22M1P U62 ( .A(n198), .B(n80), .C(n79), .D(n199), .Z(n306) );
  N1M1P U63 ( .A(n303), .Z(n199) );
  N1M1P U64 ( .A(n305), .Z(n198) );
  AOI22M1P U65 ( .A(n204), .B(n80), .C(n79), .D(n205), .Z(n294) );
  N1M1P U66 ( .A(n293), .Z(n204) );
  N1M1P U67 ( .A(n351), .Z(n153) );
  AOI22M1P U68 ( .A(n205), .B(n80), .C(n79), .D(n206), .Z(n292) );
  N1M1P U69 ( .A(n289), .Z(n206) );
  N1M1P U70 ( .A(n291), .Z(n205) );
  AOI22M1P U71 ( .A(n157), .B(n80), .C(n79), .D(n190), .Z(n324) );
  AOI22M1P U72 ( .A(n156), .B(n80), .C(n79), .D(n157), .Z(n326) );
  N1M1P U73 ( .A(n323), .Z(n157) );
  N1M1P U74 ( .A(n325), .Z(n156) );
  AOI22M1P U75 ( .A(n190), .B(n80), .C(n79), .D(n191), .Z(n322) );
  N1M1P U76 ( .A(n319), .Z(n191) );
  N1M1P U77 ( .A(n321), .Z(n190) );
  AOI22M1P U78 ( .A(n192), .B(n80), .C(n79), .D(n193), .Z(n318) );
  N1M1P U79 ( .A(n315), .Z(n193) );
  N1M1P U80 ( .A(n317), .Z(n192) );
  AOI22M1P U81 ( .A(n154), .B(n80), .C(n79), .D(n155), .Z(n330) );
  N1M1P U82 ( .A(n327), .Z(n155) );
  N1M1P U83 ( .A(n329), .Z(n154) );
  N1M1P U84 ( .A(receivedCounter[4]), .Z(n216) );
  ND2BNM1P U85 ( .B(n228), .A(n115), .Z(n86) );
  N1M1P U86 ( .A(receivedCounter[0]), .Z(n215) );
  N1M1P U87 ( .A(receivedCounter[2]), .Z(n218) );
  MUX21LM1P U88 ( .A(n345), .B(n146), .S(n75), .Z(n277) );
  N1M1P U89 ( .A(RxData[27]), .Z(n146) );
  MUX21LM1P U90 ( .A(n347), .B(n147), .S(n77), .Z(n278) );
  N1M1P U91 ( .A(RxData[28]), .Z(n147) );
  MUX21LM1P U92 ( .A(n335), .B(n141), .S(n77), .Z(n272) );
  N1M1P U93 ( .A(RxData[22]), .Z(n141) );
  MUX21LM1P U94 ( .A(n339), .B(n143), .S(n75), .Z(n274) );
  N1M1P U95 ( .A(RxData[24]), .Z(n143) );
  MUX21LM1P U96 ( .A(n353), .B(n151), .S(n75), .Z(n281) );
  N1M1P U97 ( .A(RxData[31]), .Z(n151) );
  MUX21LM1P U98 ( .A(n349), .B(n148), .S(n75), .Z(n279) );
  N1M1P U99 ( .A(RxData[29]), .Z(n148) );
  MUX21LM1P U100 ( .A(n343), .B(n145), .S(n77), .Z(n276) );
  N1M1P U101 ( .A(RxData[26]), .Z(n145) );
  MUX21LM1P U102 ( .A(n337), .B(n142), .S(n75), .Z(n273) );
  N1M1P U103 ( .A(RxData[23]), .Z(n142) );
  MUX21LM1P U104 ( .A(n351), .B(n149), .S(n75), .Z(n280) );
  N1M1P U105 ( .A(RxData[30]), .Z(n149) );
  MUX21LM1P U106 ( .A(n341), .B(n144), .S(n75), .Z(n275) );
  N1M1P U107 ( .A(RxData[25]), .Z(n144) );
  MUX21LM1P U108 ( .A(n317), .B(n132), .S(n77), .Z(n263) );
  N1M1P U109 ( .A(RxData[13]), .Z(n132) );
  MUX21LM1P U110 ( .A(n297), .B(n122), .S(n75), .Z(n253) );
  N1M1P U111 ( .A(RxData[3]), .Z(n122) );
  MUX21LM1P U112 ( .A(n323), .B(n135), .S(n77), .Z(n266) );
  N1M1P U113 ( .A(RxData[16]), .Z(n135) );
  MUX21LM1P U114 ( .A(n307), .B(n127), .S(n75), .Z(n258) );
  N1M1P U115 ( .A(RxData[8]), .Z(n127) );
  MUX21LM1P U116 ( .A(n319), .B(n133), .S(n75), .Z(n264) );
  N1M1P U117 ( .A(RxData[14]), .Z(n133) );
  MUX21LM1P U118 ( .A(n329), .B(n138), .S(n75), .Z(n269) );
  N1M1P U119 ( .A(RxData[19]), .Z(n138) );
  MUX21LM1P U120 ( .A(n293), .B(n120), .S(n75), .Z(n251) );
  N1M1P U121 ( .A(RxData[1]), .Z(n120) );
  MUX21LM1P U122 ( .A(n311), .B(n129), .S(n77), .Z(n260) );
  N1M1P U123 ( .A(RxData[10]), .Z(n129) );
  MUX21LM1P U124 ( .A(n333), .B(n140), .S(n75), .Z(n271) );
  N1M1P U125 ( .A(RxData[21]), .Z(n140) );
  MUX21LM1P U126 ( .A(n325), .B(n136), .S(n77), .Z(n267) );
  N1M1P U127 ( .A(RxData[17]), .Z(n136) );
  MUX21LM1P U128 ( .A(n291), .B(n119), .S(n75), .Z(n250) );
  N1M1P U129 ( .A(RxData[0]), .Z(n119) );
  MUX21LM1P U130 ( .A(n299), .B(n123), .S(n75), .Z(n254) );
  N1M1P U131 ( .A(RxData[4]), .Z(n123) );
  MUX21LM1P U132 ( .A(n301), .B(n124), .S(n75), .Z(n255) );
  N1M1P U133 ( .A(RxData[5]), .Z(n124) );
  MUX21LM1P U134 ( .A(n295), .B(n121), .S(n77), .Z(n252) );
  N1M1P U135 ( .A(RxData[2]), .Z(n121) );
  MUX21LM1P U136 ( .A(n321), .B(n134), .S(n75), .Z(n265) );
  N1M1P U137 ( .A(RxData[15]), .Z(n134) );
  MUX21LM1P U138 ( .A(n331), .B(n139), .S(n75), .Z(n270) );
  N1M1P U139 ( .A(RxData[20]), .Z(n139) );
  MUX21LM1P U140 ( .A(n315), .B(n131), .S(n75), .Z(n262) );
  N1M1P U141 ( .A(RxData[12]), .Z(n131) );
  MUX21LM1P U142 ( .A(n309), .B(n128), .S(n77), .Z(n259) );
  N1M1P U143 ( .A(RxData[9]), .Z(n128) );
  MUX21LM1P U144 ( .A(n303), .B(n125), .S(n75), .Z(n256) );
  N1M1P U145 ( .A(RxData[6]), .Z(n125) );
  MUX21LM1P U146 ( .A(n313), .B(n130), .S(n77), .Z(n261) );
  N1M1P U147 ( .A(RxData[11]), .Z(n130) );
  MUX21LM1P U148 ( .A(n305), .B(n126), .S(n75), .Z(n257) );
  N1M1P U149 ( .A(RxData[7]), .Z(n126) );
  MUX21LM1P U150 ( .A(n327), .B(n137), .S(n77), .Z(n268) );
  NR2M1P U151 ( .A(receivedCounter[2]), .B(receivedCounter[4]), .Z(n83) );
  ENFM1P U152 ( .A(n111), .B(n110), .Z(n112) );
  EOFM1P U153 ( .A(n109), .B(n108), .Z(n110) );
  EOFM1P U154 ( .A(n220), .B(n107), .Z(n108) );
  EOFM1P U155 ( .A(n325), .B(n106), .Z(n107) );
  ENFM1P U156 ( .A(n333), .B(n337), .Z(n106) );
  AOI22M1P U157 ( .A(n349), .B(n347), .C(n245), .D(n246), .Z(n220) );
  EOFM1P U158 ( .A(n105), .B(n219), .Z(n109) );
  AOI22M1P U159 ( .A(n345), .B(n343), .C(n243), .D(n244), .Z(n219) );
  EOFM1P U160 ( .A(n329), .B(n327), .Z(n105) );
  ENFM1P U161 ( .A(n104), .B(n103), .Z(n111) );
  ENFM1P U162 ( .A(n102), .B(n101), .Z(n103) );
  ENFM1P U163 ( .A(n323), .B(n321), .Z(n101) );
  ENFM1P U164 ( .A(n319), .B(n301), .Z(n102) );
  ENFM1P U165 ( .A(n100), .B(n99), .Z(n113) );
  ENFM1P U166 ( .A(n98), .B(n97), .Z(n99) );
  ENFM1P U167 ( .A(n96), .B(n95), .Z(n97) );
  EOFM1P U168 ( .A(n307), .B(n305), .Z(n95) );
  ENFM1P U169 ( .A(n297), .B(n303), .Z(n96) );
  ENFM1P U170 ( .A(n94), .B(n93), .Z(n98) );
  EOFM1P U171 ( .A(n293), .B(n351), .Z(n93) );
  ENFM1P U172 ( .A(n291), .B(n295), .Z(n94) );
  ENFM1P U173 ( .A(n92), .B(n91), .Z(n100) );
  ENFM1P U174 ( .A(n90), .B(n89), .Z(n91) );
  ENFM1P U175 ( .A(n317), .B(n315), .Z(n89) );
  ENFM1P U176 ( .A(n353), .B(n289), .Z(n90) );
  ENFM1P U177 ( .A(n88), .B(n87), .Z(n92) );
  ENFM1P U178 ( .A(n339), .B(n331), .Z(n87) );
  EOFM1P U179 ( .A(n335), .B(n341), .Z(n88) );
  N1M1P U180 ( .A(RxData[18]), .Z(n137) );
  N1M2P U181 ( .A(n247), .Z(n82) );
  OAI21M1P U182 ( .A(n226), .B(n227), .C(n86), .Z(n247) );
  OA21M1P U183 ( .A(n152), .B(bufferFull), .C(Core_Rcv_Ready), .Z(N243) );
  ND2M1P U184 ( .A(zeroCounter[1]), .B(zeroCounter[0]), .Z(n222) );
  NR3M1P U185 ( .A(S_Data), .B(zeroCounter[2]), .C(n222), .Z(N26) );
  N1M1P U186 ( .A(receivedCounter[5]), .Z(n240) );
  AND2M1P U187 ( .A(N26), .B(n240), .Z(N22) );
  NR3M1P U188 ( .A(S_Data), .B(zeroCounter[2]), .C(zeroCounter[0]), .Z(N24) );
  NR2BNM1P U189 ( .B(RxData_Valid), .A(Core_Rcv_Ready), .Z(n221) );
  OAI21M1P U190 ( .A(zeroCounter[1]), .B(zeroCounter[0]), .C(n222), .Z(n225)
         );
  NR3M1P U191 ( .A(S_Data), .B(zeroCounter[2]), .C(n225), .Z(N25) );
  NR2BNM1P U192 ( .B(n287), .A(dataRx), .Z(N27) );
  ND2M1P U193 ( .A(n287), .B(n78), .Z(n242) );
  N1M1P U194 ( .A(bitStuff), .Z(n227) );
  ND2BNM1P U195 ( .B(n242), .A(n82), .Z(n248) );
  ND2M1P U196 ( .A(n79), .B(n215), .Z(n229) );
  OAI211M1P U197 ( .A(n82), .B(n215), .C(n287), .D(n229), .Z(n249) );
  AOI21M1P U198 ( .A(n79), .B(n215), .C(n81), .Z(n230) );
  N1M1P U199 ( .A(receivedCounter[1]), .Z(n234) );
  NR2M1P U200 ( .A(receivedCounter[1]), .B(n78), .Z(n231) );
  OAI22CDNM1P U201 ( .A(n230), .B(n234), .C(receivedCounter[0]), .D(n231), .Z(
        n282) );
  AOI211M1P U202 ( .A(n79), .B(n215), .C(n231), .D(n81), .Z(n233) );
  ND3M1P U203 ( .A(receivedCounter[1]), .B(receivedCounter[0]), .C(n79), .Z(
        n232) );
  AOI22M1P U204 ( .A(receivedCounter[2]), .B(n233), .C(n232), .D(n218), .Z(
        n283) );
  NR3M1P U205 ( .A(n234), .B(n218), .C(n215), .Z(n238) );
  N1M1P U206 ( .A(n238), .Z(n235) );
  AOI21M1P U207 ( .A(n235), .B(n79), .C(n81), .Z(n237) );
  ND2M1P U208 ( .A(n79), .B(n217), .Z(n236) );
  OAI22M1P U209 ( .A(n237), .B(n217), .C(n236), .D(n235), .Z(n284) );
  OA21M1P U210 ( .A(n78), .B(receivedCounter[3]), .C(n237), .Z(n241) );
  ND3M1P U211 ( .A(receivedCounter[3]), .B(n79), .C(n238), .Z(n239) );
  AOI22M1P U212 ( .A(receivedCounter[4]), .B(n241), .C(n239), .D(n216), .Z(
        n285) );
  OAI22M1P U213 ( .A(n241), .B(n240), .C(n216), .D(n239), .Z(n286) );
  ND2BNM1P U214 ( .B(S_Data), .A(zeroCounter[2]), .Z(n288) );
  AOI22M1P U215 ( .A(n79), .B(n209), .C(n210), .D(n81), .Z(n334) );
  AOI22M1P U216 ( .A(n79), .B(n210), .C(n211), .D(n81), .Z(n336) );
  AOI22M1P U217 ( .A(n79), .B(n211), .C(n212), .D(n81), .Z(n338) );
  AOI22M1P U218 ( .A(n79), .B(n212), .C(n213), .D(n81), .Z(n340) );
  AOI22M1P U219 ( .A(n79), .B(n213), .C(n214), .D(n81), .Z(n342) );
  AOI22M1P U220 ( .A(n79), .B(n214), .C(n243), .D(n81), .Z(n344) );
  AOI22M1P U221 ( .A(n79), .B(n243), .C(n244), .D(n81), .Z(n346) );
  AOI22M1P U222 ( .A(n79), .B(n244), .C(n245), .D(n81), .Z(n348) );
  AOI22M1P U223 ( .A(n79), .B(n245), .C(n246), .D(n81), .Z(n350) );
endmodule


module rx_2 ( Clk_s, Rst_n, Core_Rcv_Ready, S_Data, RxData_Valid, RxData, 
        Rx_Ready, Rx_Error );
  output [31:0] RxData;
  input Clk_s, Rst_n, Core_Rcv_Ready, S_Data;
  output RxData_Valid, Rx_Ready, Rx_Error;
  wire   bitStuff, N22, N24, N25, N26, dataRx, bufferFull, N27, N229, N242,
         N243, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352;
  wire   [2:0] zeroCounter;
  wire   [5:0] receivedCounter;

  FD4QM1P startSeq_reg ( .D(n286), .CP(Clk_s), .SD(Rst_n), .Q(n285) );
  FD2QM1P \receivedCounter_reg[5]  ( .D(n284), .CP(Clk_s), .CD(Rst_n), .Q(
        receivedCounter[5]) );
  FD4QM1P \receivedPacket_reg[0]  ( .D(n288), .CP(Clk_s), .SD(Rst_n), .Q(n287)
         );
  FD4QM1P \receivedPacket_reg[1]  ( .D(n290), .CP(Clk_s), .SD(Rst_n), .Q(n289)
         );
  FD4QM1P \receivedPacket_reg[2]  ( .D(n292), .CP(Clk_s), .SD(Rst_n), .Q(n291)
         );
  FD4QM1P \receivedPacket_reg[3]  ( .D(n294), .CP(Clk_s), .SD(Rst_n), .Q(n293)
         );
  FD4QM1P \receivedPacket_reg[4]  ( .D(n296), .CP(Clk_s), .SD(Rst_n), .Q(n295)
         );
  FD4QM1P \receivedPacket_reg[5]  ( .D(n298), .CP(Clk_s), .SD(Rst_n), .Q(n297)
         );
  FD4QM1P \receivedPacket_reg[6]  ( .D(n300), .CP(Clk_s), .SD(Rst_n), .Q(n299)
         );
  FD4QM1P \receivedPacket_reg[7]  ( .D(n302), .CP(Clk_s), .SD(Rst_n), .Q(n301)
         );
  FD4QM1P \receivedPacket_reg[8]  ( .D(n304), .CP(Clk_s), .SD(Rst_n), .Q(n303)
         );
  FD4QM1P \receivedPacket_reg[9]  ( .D(n306), .CP(Clk_s), .SD(Rst_n), .Q(n305)
         );
  FD4QM1P \receivedPacket_reg[10]  ( .D(n308), .CP(Clk_s), .SD(Rst_n), .Q(n307) );
  FD4QM1P \receivedPacket_reg[11]  ( .D(n310), .CP(Clk_s), .SD(Rst_n), .Q(n309) );
  FD4QM1P \receivedPacket_reg[12]  ( .D(n312), .CP(Clk_s), .SD(Rst_n), .Q(n311) );
  FD4QM1P \receivedPacket_reg[13]  ( .D(n314), .CP(Clk_s), .SD(Rst_n), .Q(n313) );
  FD4QM1P \receivedPacket_reg[14]  ( .D(n316), .CP(Clk_s), .SD(Rst_n), .Q(n315) );
  FD4QM1P \receivedPacket_reg[15]  ( .D(n318), .CP(Clk_s), .SD(Rst_n), .Q(n317) );
  FD4QM1P \receivedPacket_reg[16]  ( .D(n320), .CP(Clk_s), .SD(Rst_n), .Q(n319) );
  FD4QM1P \receivedPacket_reg[17]  ( .D(n322), .CP(Clk_s), .SD(Rst_n), .Q(n321) );
  FD4QM1P \receivedPacket_reg[18]  ( .D(n324), .CP(Clk_s), .SD(Rst_n), .Q(n323) );
  FD4QM1P \receivedPacket_reg[19]  ( .D(n326), .CP(Clk_s), .SD(Rst_n), .Q(n325) );
  FD4QM1P \receivedPacket_reg[20]  ( .D(n328), .CP(Clk_s), .SD(Rst_n), .Q(n327) );
  FD4QM1P \receivedPacket_reg[21]  ( .D(n330), .CP(Clk_s), .SD(Rst_n), .Q(n329) );
  FD4QM1P \receivedPacket_reg[23]  ( .D(n334), .CP(Clk_s), .SD(Rst_n), .Q(n333) );
  FD4QM1P \receivedPacket_reg[25]  ( .D(n338), .CP(Clk_s), .SD(Rst_n), .Q(n337) );
  FD4QM1P \receivedPacket_reg[26]  ( .D(n340), .CP(Clk_s), .SD(Rst_n), .Q(n339) );
  FD4QM1P \receivedPacket_reg[29]  ( .D(n346), .CP(Clk_s), .SD(Rst_n), .Q(n345) );
  FD4QM1P \receivedPacket_reg[31]  ( .D(n350), .CP(Clk_s), .SD(Rst_n), .Q(n349) );
  FD4QM1P \receivedPacket_reg[32]  ( .D(n352), .CP(Clk_s), .SD(Rst_n), .Q(n351) );
  FD2QM1P \RxData_reg[31]  ( .D(n279), .CP(Clk_s), .CD(Rst_n), .Q(RxData[31])
         );
  FD2QM1P \RxData_reg[30]  ( .D(n278), .CP(Clk_s), .CD(Rst_n), .Q(RxData[30])
         );
  FD2QM1P \RxData_reg[29]  ( .D(n277), .CP(Clk_s), .CD(Rst_n), .Q(RxData[29])
         );
  FD2QM1P \RxData_reg[28]  ( .D(n276), .CP(Clk_s), .CD(Rst_n), .Q(RxData[28])
         );
  FD2QM1P \RxData_reg[27]  ( .D(n275), .CP(Clk_s), .CD(Rst_n), .Q(RxData[27])
         );
  FD2QM1P \RxData_reg[26]  ( .D(n274), .CP(Clk_s), .CD(Rst_n), .Q(RxData[26])
         );
  FD2QM1P \RxData_reg[25]  ( .D(n273), .CP(Clk_s), .CD(Rst_n), .Q(RxData[25])
         );
  FD2QM1P \RxData_reg[24]  ( .D(n272), .CP(Clk_s), .CD(Rst_n), .Q(RxData[24])
         );
  FD2QM1P \RxData_reg[23]  ( .D(n271), .CP(Clk_s), .CD(Rst_n), .Q(RxData[23])
         );
  FD2QM1P \RxData_reg[22]  ( .D(n270), .CP(Clk_s), .CD(Rst_n), .Q(RxData[22])
         );
  FD2QM1P \RxData_reg[21]  ( .D(n269), .CP(Clk_s), .CD(Rst_n), .Q(RxData[21])
         );
  FD2QM1P \RxData_reg[20]  ( .D(n268), .CP(Clk_s), .CD(Rst_n), .Q(RxData[20])
         );
  FD2QM1P \RxData_reg[19]  ( .D(n267), .CP(Clk_s), .CD(Rst_n), .Q(RxData[19])
         );
  FD2QM1P \RxData_reg[18]  ( .D(n266), .CP(Clk_s), .CD(Rst_n), .Q(RxData[18])
         );
  FD2QM1P \RxData_reg[17]  ( .D(n265), .CP(Clk_s), .CD(Rst_n), .Q(RxData[17])
         );
  FD2QM1P \RxData_reg[16]  ( .D(n264), .CP(Clk_s), .CD(Rst_n), .Q(RxData[16])
         );
  FD2QM1P \RxData_reg[15]  ( .D(n263), .CP(Clk_s), .CD(Rst_n), .Q(RxData[15])
         );
  FD2QM1P \RxData_reg[14]  ( .D(n262), .CP(Clk_s), .CD(Rst_n), .Q(RxData[14])
         );
  FD2QM1P \RxData_reg[13]  ( .D(n261), .CP(Clk_s), .CD(Rst_n), .Q(RxData[13])
         );
  FD2QM1P \RxData_reg[12]  ( .D(n260), .CP(Clk_s), .CD(Rst_n), .Q(RxData[12])
         );
  FD2QM1P \RxData_reg[11]  ( .D(n259), .CP(Clk_s), .CD(Rst_n), .Q(RxData[11])
         );
  FD2QM1P \RxData_reg[10]  ( .D(n258), .CP(Clk_s), .CD(Rst_n), .Q(RxData[10])
         );
  FD2QM1P \RxData_reg[9]  ( .D(n257), .CP(Clk_s), .CD(Rst_n), .Q(RxData[9]) );
  FD2QM1P \RxData_reg[8]  ( .D(n256), .CP(Clk_s), .CD(Rst_n), .Q(RxData[8]) );
  FD2QM1P \RxData_reg[7]  ( .D(n255), .CP(Clk_s), .CD(Rst_n), .Q(RxData[7]) );
  FD2QM1P \RxData_reg[6]  ( .D(n254), .CP(Clk_s), .CD(Rst_n), .Q(RxData[6]) );
  FD2QM1P \RxData_reg[5]  ( .D(n253), .CP(Clk_s), .CD(Rst_n), .Q(RxData[5]) );
  FD2QM1P \RxData_reg[4]  ( .D(n252), .CP(Clk_s), .CD(Rst_n), .Q(RxData[4]) );
  FD2QM1P \RxData_reg[3]  ( .D(n251), .CP(Clk_s), .CD(Rst_n), .Q(RxData[3]) );
  FD2QM1P \RxData_reg[2]  ( .D(n250), .CP(Clk_s), .CD(Rst_n), .Q(RxData[2]) );
  FD2QM1P \RxData_reg[1]  ( .D(n249), .CP(Clk_s), .CD(Rst_n), .Q(RxData[1]) );
  FD2QM1P \RxData_reg[0]  ( .D(n248), .CP(Clk_s), .CD(Rst_n), .Q(RxData[0]) );
  FD2QM1P \receivedCounter_reg[4]  ( .D(n283), .CP(Clk_s), .CD(Rst_n), .Q(
        receivedCounter[4]) );
  FD4QM1P \receivedPacket_reg[24]  ( .D(n336), .CP(Clk_s), .SD(Rst_n), .Q(n335) );
  FD4QM3P \receivedPacket_reg[28]  ( .D(n344), .CP(Clk_s), .SD(Rst_n), .Q(n343) );
  FD4QM3P \receivedPacket_reg[22]  ( .D(n332), .CP(Clk_s), .SD(Rst_n), .Q(n331) );
  FD4QM3P \receivedPacket_reg[30]  ( .D(n348), .CP(Clk_s), .SD(Rst_n), .Q(n347) );
  FD4QM3P \receivedPacket_reg[27]  ( .D(n342), .CP(Clk_s), .SD(Rst_n), .Q(n341) );
  FD2QM1P \zeroCounter_reg[0]  ( .D(N24), .CP(Clk_s), .CD(Rst_n), .Q(
        zeroCounter[0]) );
  FD2QM1P Rx_Ready_reg ( .D(N27), .CP(Clk_s), .CD(Rst_n), .Q(Rx_Ready) );
  FD2QM1P \zeroCounter_reg[1]  ( .D(N25), .CP(Clk_s), .CD(Rst_n), .Q(
        zeroCounter[1]) );
  FD2QM1P \zeroCounter_reg[2]  ( .D(N26), .CP(Clk_s), .CD(Rst_n), .Q(
        zeroCounter[2]) );
  FD2QM1P bitStuff_reg ( .D(N22), .CP(Clk_s), .CD(Rst_n), .Q(bitStuff) );
  FD2QM1P dataRx_reg ( .D(n246), .CP(Clk_s), .CD(Rst_n), .Q(dataRx) );
  FD2QM1P Rx_Error_reg ( .D(N229), .CP(Clk_s), .CD(Rst_n), .Q(Rx_Error) );
  FD2QM1P \receivedCounter_reg[0]  ( .D(n247), .CP(Clk_s), .CD(Rst_n), .Q(
        receivedCounter[0]) );
  FD2QM1P bufferFull_reg ( .D(N242), .CP(Clk_s), .CD(Rst_n), .Q(bufferFull) );
  FD2QM1P \receivedCounter_reg[1]  ( .D(n280), .CP(Clk_s), .CD(Rst_n), .Q(
        receivedCounter[1]) );
  FD2QM1P RxData_Valid_reg ( .D(N243), .CP(Clk_s), .CD(Rst_n), .Q(RxData_Valid) );
  FD2QM1P \receivedCounter_reg[3]  ( .D(n282), .CP(Clk_s), .CD(Rst_n), .Q(
        receivedCounter[3]) );
  FD2QM1P \receivedCounter_reg[2]  ( .D(n281), .CP(Clk_s), .CD(Rst_n), .Q(
        receivedCounter[2]) );
  ND2M1P U3 ( .A(dataRx), .B(n285), .Z(n222) );
  ND2M1P U4 ( .A(n116), .B(n114), .Z(n74) );
  NR2BNM1P U5 ( .B(n116), .A(n114), .Z(n113) );
  N1M1P U6 ( .A(n341), .Z(n241) );
  N1M1P U7 ( .A(n347), .Z(n244) );
  N1M1P U8 ( .A(n343), .Z(n242) );
  N1M3P U9 ( .A(n74), .Z(n75) );
  N1M2P U10 ( .A(n78), .Z(n76) );
  AOI22DNM1P U11 ( .A(n151), .B(n75), .D(n351), .C(n76), .Z(n352) );
  ND2FM3P U12 ( .A(n112), .B(n226), .Z(n115) );
  ND2M10P U13 ( .A(n205), .B(n116), .Z(n148) );
  NR2M6P U14 ( .A(n115), .B(n114), .Z(n205) );
  N1M2P U15 ( .A(n345), .Z(n243) );
  AOI22M2P U16 ( .A(n343), .B(n341), .C(n241), .D(n242), .Z(n217) );
  ENM2P U17 ( .A(n111), .B(n110), .Z(n112) );
  N1M3P U18 ( .A(n78), .Z(n77) );
  NR2FM1P U19 ( .A(n222), .B(bitStuff), .Z(n116) );
  OAI21M2P U20 ( .A(n81), .B(n80), .C(receivedCounter[5]), .Z(n114) );
  N1M1P U21 ( .A(bufferFull), .Z(n226) );
  OR2M1P U22 ( .A(receivedCounter[3]), .B(receivedCounter[0]), .Z(n80) );
  ND2BNM1P U23 ( .B(receivedCounter[1]), .A(n79), .Z(n81) );
  AOI22M1P U24 ( .A(n151), .B(n77), .C(n244), .D(n75), .Z(n350) );
  N1M1P U25 ( .A(n337), .Z(n211) );
  N1M1P U26 ( .A(n339), .Z(n212) );
  N1M1P U27 ( .A(n331), .Z(n208) );
  N1M1P U28 ( .A(n335), .Z(n210) );
  N1M1P U29 ( .A(n333), .Z(n209) );
  AOI22M1P U30 ( .A(n207), .B(n77), .C(n75), .D(n152), .Z(n330) );
  N1M1P U31 ( .A(n329), .Z(n207) );
  OAI21M1P U32 ( .A(n226), .B(n219), .C(n206), .Z(N242) );
  N1M1P U33 ( .A(receivedCounter[3]), .Z(n215) );
  AOI22M1P U34 ( .A(n204), .B(n76), .C(n240), .D(S_Data), .Z(n288) );
  N1M1P U35 ( .A(receivedCounter[4]), .Z(n214) );
  N1M1P U36 ( .A(receivedCounter[0]), .Z(n213) );
  N1M1P U37 ( .A(receivedCounter[2]), .Z(n216) );
  AOI22M1P U38 ( .A(n201), .B(n76), .C(n75), .D(n202), .Z(n294) );
  AOI22M1P U39 ( .A(n203), .B(n76), .C(n75), .D(n204), .Z(n290) );
  N1M1P U40 ( .A(n287), .Z(n204) );
  AOI22M1P U41 ( .A(n153), .B(n76), .C(n75), .D(n154), .Z(n326) );
  AOI22M1P U42 ( .A(n152), .B(n76), .C(n75), .D(n153), .Z(n328) );
  N1M1P U43 ( .A(n325), .Z(n153) );
  N1M1P U44 ( .A(n327), .Z(n152) );
  AOI22M1P U45 ( .A(n199), .B(n76), .C(n75), .D(n200), .Z(n298) );
  AOI22M1P U46 ( .A(n155), .B(n76), .C(n75), .D(n156), .Z(n322) );
  AOI22M1P U47 ( .A(n198), .B(n76), .C(n75), .D(n199), .Z(n300) );
  N1M1P U48 ( .A(n297), .Z(n199) );
  AOI22M1P U49 ( .A(n200), .B(n76), .C(n75), .D(n201), .Z(n296) );
  N1M1P U50 ( .A(n293), .Z(n201) );
  N1M1P U51 ( .A(n295), .Z(n200) );
  AOI22M1P U52 ( .A(n202), .B(n76), .C(n75), .D(n203), .Z(n292) );
  N1M1P U53 ( .A(n289), .Z(n203) );
  N1M1P U54 ( .A(n291), .Z(n202) );
  N1M1P U55 ( .A(n349), .Z(n151) );
  AOI22M1P U56 ( .A(n197), .B(n76), .C(n75), .D(n198), .Z(n302) );
  N1M1P U57 ( .A(n299), .Z(n198) );
  AOI22M1P U58 ( .A(n156), .B(n76), .C(n75), .D(n157), .Z(n320) );
  N1M1P U59 ( .A(n319), .Z(n156) );
  AOI22M1P U60 ( .A(n154), .B(n76), .C(n75), .D(n155), .Z(n324) );
  N1M1P U61 ( .A(n321), .Z(n155) );
  N1M1P U62 ( .A(n323), .Z(n154) );
  AOI22M1P U63 ( .A(n196), .B(n76), .C(n75), .D(n197), .Z(n304) );
  N1M1P U64 ( .A(n301), .Z(n197) );
  AOI22M1P U65 ( .A(n192), .B(n76), .C(n75), .D(n193), .Z(n312) );
  AOI22M1P U66 ( .A(n195), .B(n76), .C(n75), .D(n196), .Z(n306) );
  N1M1P U67 ( .A(n303), .Z(n196) );
  AOI22M1P U68 ( .A(n194), .B(n76), .C(n75), .D(n195), .Z(n308) );
  N1M1P U69 ( .A(n305), .Z(n195) );
  AOI22M1P U70 ( .A(n193), .B(n76), .C(n75), .D(n194), .Z(n310) );
  N1M1P U71 ( .A(n307), .Z(n194) );
  N1M1P U72 ( .A(n309), .Z(n193) );
  AOI22M1P U73 ( .A(n190), .B(n76), .C(n75), .D(n191), .Z(n316) );
  AOI22M1P U74 ( .A(n157), .B(n76), .C(n75), .D(n190), .Z(n318) );
  N1M1P U75 ( .A(n315), .Z(n190) );
  N1M1P U76 ( .A(n317), .Z(n157) );
  AOI22M1P U77 ( .A(n191), .B(n76), .C(n75), .D(n192), .Z(n314) );
  N1M1P U78 ( .A(n311), .Z(n192) );
  ND2BNM1P U79 ( .B(n226), .A(n113), .Z(n82) );
  N1M1P U80 ( .A(n313), .Z(n191) );
  MUX21LM1P U81 ( .A(n343), .B(n144), .S(n148), .Z(n275) );
  N1M1P U82 ( .A(RxData[27]), .Z(n144) );
  MUX21LM1P U83 ( .A(n341), .B(n143), .S(n148), .Z(n274) );
  N1M1P U84 ( .A(RxData[26]), .Z(n143) );
  MUX21LM1P U85 ( .A(n345), .B(n145), .S(n148), .Z(n276) );
  N1M1P U86 ( .A(RxData[28]), .Z(n145) );
  MUX21LM1P U87 ( .A(n347), .B(n146), .S(n148), .Z(n277) );
  N1M1P U88 ( .A(RxData[29]), .Z(n146) );
  MUX21LM1P U89 ( .A(n333), .B(n139), .S(n148), .Z(n270) );
  N1M1P U90 ( .A(RxData[22]), .Z(n139) );
  MUX21LM1P U91 ( .A(n351), .B(n149), .S(n148), .Z(n279) );
  N1M1P U92 ( .A(RxData[31]), .Z(n149) );
  MUX21LM1P U93 ( .A(n337), .B(n141), .S(n148), .Z(n272) );
  N1M1P U94 ( .A(RxData[24]), .Z(n141) );
  MUX21LM1P U95 ( .A(n339), .B(n142), .S(n148), .Z(n273) );
  N1M1P U96 ( .A(RxData[25]), .Z(n142) );
  MUX21LM1P U97 ( .A(n349), .B(n147), .S(n148), .Z(n278) );
  N1M1P U98 ( .A(RxData[30]), .Z(n147) );
  MUX21LM1P U99 ( .A(n335), .B(n140), .S(n148), .Z(n271) );
  N1M1P U100 ( .A(RxData[23]), .Z(n140) );
  MUX21LM1P U101 ( .A(n317), .B(n131), .S(n148), .Z(n262) );
  N1M1P U102 ( .A(RxData[14]), .Z(n131) );
  MUX21LM1P U103 ( .A(n297), .B(n121), .S(n148), .Z(n252) );
  N1M1P U104 ( .A(RxData[4]), .Z(n121) );
  MUX21LM1P U105 ( .A(n309), .B(n127), .S(n148), .Z(n258) );
  N1M1P U106 ( .A(RxData[10]), .Z(n127) );
  MUX21LM1P U107 ( .A(n327), .B(n136), .S(n148), .Z(n267) );
  N1M1P U108 ( .A(RxData[19]), .Z(n136) );
  MUX21LM1P U109 ( .A(n321), .B(n133), .S(n148), .Z(n264) );
  N1M1P U110 ( .A(RxData[16]), .Z(n133) );
  MUX21LM1P U111 ( .A(n291), .B(n118), .S(n148), .Z(n249) );
  N1M1P U112 ( .A(RxData[1]), .Z(n118) );
  MUX21LM1P U113 ( .A(n289), .B(n117), .S(n148), .Z(n248) );
  N1M1P U114 ( .A(RxData[0]), .Z(n117) );
  MUX21LM1P U115 ( .A(n305), .B(n125), .S(n148), .Z(n256) );
  N1M1P U116 ( .A(RxData[8]), .Z(n125) );
  MUX21LM1P U117 ( .A(n323), .B(n134), .S(n148), .Z(n265) );
  N1M1P U118 ( .A(RxData[17]), .Z(n134) );
  MUX21LM1P U119 ( .A(n315), .B(n130), .S(n148), .Z(n261) );
  N1M1P U120 ( .A(RxData[13]), .Z(n130) );
  MUX21LM1P U121 ( .A(n295), .B(n120), .S(n148), .Z(n251) );
  N1M1P U122 ( .A(RxData[3]), .Z(n120) );
  MUX21LM1P U123 ( .A(n313), .B(n129), .S(n148), .Z(n260) );
  N1M1P U124 ( .A(RxData[12]), .Z(n129) );
  MUX21LM1P U125 ( .A(n301), .B(n123), .S(n148), .Z(n254) );
  N1M1P U126 ( .A(RxData[6]), .Z(n123) );
  MUX21LM1P U127 ( .A(n319), .B(n132), .S(n148), .Z(n263) );
  N1M1P U128 ( .A(RxData[15]), .Z(n132) );
  MUX21LM1P U129 ( .A(n293), .B(n119), .S(n148), .Z(n250) );
  N1M1P U130 ( .A(RxData[2]), .Z(n119) );
  MUX21LM1P U131 ( .A(n307), .B(n126), .S(n148), .Z(n257) );
  N1M1P U132 ( .A(RxData[9]), .Z(n126) );
  MUX21LM1P U133 ( .A(n299), .B(n122), .S(n148), .Z(n253) );
  N1M1P U134 ( .A(RxData[5]), .Z(n122) );
  MUX21LM1P U135 ( .A(n329), .B(n137), .S(n148), .Z(n268) );
  N1M1P U136 ( .A(RxData[20]), .Z(n137) );
  MUX21LM1P U137 ( .A(n303), .B(n124), .S(n148), .Z(n255) );
  N1M1P U138 ( .A(RxData[7]), .Z(n124) );
  MUX21LM1P U139 ( .A(n311), .B(n128), .S(n148), .Z(n259) );
  N1M1P U140 ( .A(RxData[11]), .Z(n128) );
  MUX21LM1P U141 ( .A(n325), .B(n135), .S(n148), .Z(n266) );
  N1M1P U142 ( .A(RxData[18]), .Z(n135) );
  MUX21LM1P U143 ( .A(n331), .B(n138), .S(n148), .Z(n269) );
  NR2M1P U144 ( .A(receivedCounter[2]), .B(receivedCounter[4]), .Z(n79) );
  ENFM1P U145 ( .A(n109), .B(n108), .Z(n110) );
  EOFM1P U146 ( .A(n107), .B(n106), .Z(n108) );
  EOFM1P U147 ( .A(n218), .B(n105), .Z(n106) );
  EOFM1P U148 ( .A(n323), .B(n104), .Z(n105) );
  ENFM1P U149 ( .A(n331), .B(n335), .Z(n104) );
  EOFM1P U150 ( .A(n327), .B(n325), .Z(n103) );
  ENFM1P U151 ( .A(n102), .B(n101), .Z(n109) );
  ENFM1P U152 ( .A(n100), .B(n99), .Z(n101) );
  ENFM1P U153 ( .A(n321), .B(n319), .Z(n99) );
  ENFM1P U154 ( .A(n317), .B(n299), .Z(n100) );
  ENFM1P U155 ( .A(n98), .B(n97), .Z(n102) );
  EOFM1P U156 ( .A(n297), .B(n311), .Z(n97) );
  ENFM1P U157 ( .A(n309), .B(n307), .Z(n98) );
  ENFM1P U158 ( .A(n96), .B(n95), .Z(n111) );
  ENFM1P U159 ( .A(n94), .B(n93), .Z(n95) );
  ENFM1P U160 ( .A(n92), .B(n91), .Z(n93) );
  EOFM1P U161 ( .A(n305), .B(n303), .Z(n91) );
  ENFM1P U162 ( .A(n295), .B(n301), .Z(n92) );
  ENFM1P U163 ( .A(n90), .B(n89), .Z(n94) );
  EOFM1P U164 ( .A(n291), .B(n349), .Z(n89) );
  ENFM1P U165 ( .A(n289), .B(n293), .Z(n90) );
  ENFM1P U166 ( .A(n88), .B(n87), .Z(n96) );
  ENFM1P U167 ( .A(n86), .B(n85), .Z(n87) );
  ENFM1P U168 ( .A(n315), .B(n313), .Z(n85) );
  ENFM1P U169 ( .A(n351), .B(n287), .Z(n86) );
  ENFM1P U170 ( .A(n84), .B(n83), .Z(n88) );
  ENFM1P U171 ( .A(n337), .B(n329), .Z(n83) );
  EOFM1P U172 ( .A(n333), .B(n339), .Z(n84) );
  N1M1P U173 ( .A(RxData[21]), .Z(n138) );
  N1M2P U174 ( .A(n245), .Z(n78) );
  OAI21M1P U175 ( .A(n222), .B(n225), .C(n82), .Z(n245) );
  AND3M1P U176 ( .A(n115), .B(n113), .C(n226), .Z(N229) );
  N1M1P U177 ( .A(n205), .Z(n206) );
  NR2BNM1P U178 ( .B(RxData_Valid), .A(n205), .Z(n150) );
  EOFM1P U179 ( .A(n103), .B(n217), .Z(n107) );
  OA21M1P U180 ( .A(n150), .B(bufferFull), .C(Core_Rcv_Ready), .Z(N243) );
  ND2M1P U181 ( .A(zeroCounter[1]), .B(zeroCounter[0]), .Z(n220) );
  NR3M1P U182 ( .A(S_Data), .B(zeroCounter[2]), .C(n220), .Z(N26) );
  N1M1P U183 ( .A(receivedCounter[5]), .Z(n238) );
  AND2M1P U184 ( .A(N26), .B(n238), .Z(N22) );
  AOI22M1P U185 ( .A(n347), .B(n345), .C(n243), .D(n244), .Z(n218) );
  NR3M1P U186 ( .A(S_Data), .B(zeroCounter[2]), .C(zeroCounter[0]), .Z(N24) );
  NR2BNM1P U187 ( .B(RxData_Valid), .A(Core_Rcv_Ready), .Z(n219) );
  OAI21M1P U188 ( .A(zeroCounter[1]), .B(zeroCounter[0]), .C(n220), .Z(n221)
         );
  NR3M1P U189 ( .A(S_Data), .B(zeroCounter[2]), .C(n221), .Z(N25) );
  NR2BNM1P U190 ( .B(n285), .A(dataRx), .Z(N27) );
  ND2M1P U191 ( .A(n285), .B(n74), .Z(n240) );
  N1M1P U192 ( .A(bitStuff), .Z(n225) );
  ND2BNM1P U193 ( .B(n240), .A(n78), .Z(n246) );
  ND2M1P U194 ( .A(n75), .B(n213), .Z(n227) );
  OAI211M1P U195 ( .A(n78), .B(n213), .C(n285), .D(n227), .Z(n247) );
  AOI21M1P U196 ( .A(n75), .B(n213), .C(n77), .Z(n228) );
  N1M1P U197 ( .A(receivedCounter[1]), .Z(n232) );
  NR2M1P U198 ( .A(receivedCounter[1]), .B(n74), .Z(n229) );
  OAI22CDNM1P U199 ( .A(n228), .B(n232), .C(receivedCounter[0]), .D(n229), .Z(
        n280) );
  AOI211M1P U200 ( .A(n75), .B(n213), .C(n229), .D(n77), .Z(n231) );
  ND3M1P U201 ( .A(receivedCounter[1]), .B(receivedCounter[0]), .C(n75), .Z(
        n230) );
  AOI22M1P U202 ( .A(receivedCounter[2]), .B(n231), .C(n230), .D(n216), .Z(
        n281) );
  NR3M1P U203 ( .A(n232), .B(n216), .C(n213), .Z(n236) );
  N1M1P U204 ( .A(n236), .Z(n233) );
  AOI21M1P U205 ( .A(n233), .B(n75), .C(n77), .Z(n235) );
  ND2M1P U206 ( .A(n75), .B(n215), .Z(n234) );
  OAI22M1P U207 ( .A(n235), .B(n215), .C(n234), .D(n233), .Z(n282) );
  OA21M1P U208 ( .A(n74), .B(receivedCounter[3]), .C(n235), .Z(n239) );
  ND3M1P U209 ( .A(receivedCounter[3]), .B(n75), .C(n236), .Z(n237) );
  AOI22M1P U210 ( .A(receivedCounter[4]), .B(n239), .C(n237), .D(n214), .Z(
        n283) );
  OAI22M1P U211 ( .A(n239), .B(n238), .C(n214), .D(n237), .Z(n284) );
  ND2BNM1P U212 ( .B(S_Data), .A(zeroCounter[2]), .Z(n286) );
  AOI22M1P U213 ( .A(n75), .B(n207), .C(n208), .D(n77), .Z(n332) );
  AOI22M1P U214 ( .A(n75), .B(n208), .C(n209), .D(n77), .Z(n334) );
  AOI22M1P U215 ( .A(n75), .B(n209), .C(n210), .D(n77), .Z(n336) );
  AOI22M1P U216 ( .A(n75), .B(n210), .C(n211), .D(n77), .Z(n338) );
  AOI22M1P U217 ( .A(n75), .B(n211), .C(n212), .D(n77), .Z(n340) );
  AOI22M1P U218 ( .A(n75), .B(n212), .C(n241), .D(n77), .Z(n342) );
  AOI22M1P U219 ( .A(n75), .B(n241), .C(n242), .D(n77), .Z(n344) );
  AOI22M1P U220 ( .A(n75), .B(n242), .C(n243), .D(n77), .Z(n346) );
  AOI22M1P U221 ( .A(n75), .B(n243), .C(n244), .D(n77), .Z(n348) );
endmodule


module rx_3 ( Clk_s, Rst_n, Core_Rcv_Ready, S_Data, RxData_Valid, RxData, 
        Rx_Ready, Rx_Error );
  output [31:0] RxData;
  input Clk_s, Rst_n, Core_Rcv_Ready, S_Data;
  output RxData_Valid, Rx_Ready, Rx_Error;
  wire   bitStuff, N22, N24, N25, N26, dataRx, bufferFull, N27, N229, N242,
         N243, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353;
  wire   [2:0] zeroCounter;
  wire   [5:0] receivedCounter;

  FD4QM1P startSeq_reg ( .D(n287), .CP(Clk_s), .SD(Rst_n), .Q(n286) );
  FD4QM1P \receivedPacket_reg[0]  ( .D(n289), .CP(Clk_s), .SD(Rst_n), .Q(n288)
         );
  FD4QM1P \receivedPacket_reg[1]  ( .D(n291), .CP(Clk_s), .SD(Rst_n), .Q(n290)
         );
  FD4QM1P \receivedPacket_reg[2]  ( .D(n293), .CP(Clk_s), .SD(Rst_n), .Q(n292)
         );
  FD4QM1P \receivedPacket_reg[3]  ( .D(n295), .CP(Clk_s), .SD(Rst_n), .Q(n294)
         );
  FD4QM1P \receivedPacket_reg[4]  ( .D(n297), .CP(Clk_s), .SD(Rst_n), .Q(n296)
         );
  FD4QM1P \receivedPacket_reg[5]  ( .D(n299), .CP(Clk_s), .SD(Rst_n), .Q(n298)
         );
  FD4QM1P \receivedPacket_reg[6]  ( .D(n301), .CP(Clk_s), .SD(Rst_n), .Q(n300)
         );
  FD4QM1P \receivedPacket_reg[7]  ( .D(n303), .CP(Clk_s), .SD(Rst_n), .Q(n302)
         );
  FD4QM1P \receivedPacket_reg[8]  ( .D(n305), .CP(Clk_s), .SD(Rst_n), .Q(n304)
         );
  FD4QM1P \receivedPacket_reg[9]  ( .D(n307), .CP(Clk_s), .SD(Rst_n), .Q(n306)
         );
  FD4QM1P \receivedPacket_reg[10]  ( .D(n309), .CP(Clk_s), .SD(Rst_n), .Q(n308) );
  FD4QM1P \receivedPacket_reg[11]  ( .D(n311), .CP(Clk_s), .SD(Rst_n), .Q(n310) );
  FD4QM1P \receivedPacket_reg[12]  ( .D(n313), .CP(Clk_s), .SD(Rst_n), .Q(n312) );
  FD4QM1P \receivedPacket_reg[13]  ( .D(n315), .CP(Clk_s), .SD(Rst_n), .Q(n314) );
  FD4QM1P \receivedPacket_reg[14]  ( .D(n317), .CP(Clk_s), .SD(Rst_n), .Q(n316) );
  FD4QM1P \receivedPacket_reg[15]  ( .D(n319), .CP(Clk_s), .SD(Rst_n), .Q(n318) );
  FD4QM1P \receivedPacket_reg[16]  ( .D(n321), .CP(Clk_s), .SD(Rst_n), .Q(n320) );
  FD4QM1P \receivedPacket_reg[17]  ( .D(n323), .CP(Clk_s), .SD(Rst_n), .Q(n322) );
  FD4QM1P \receivedPacket_reg[18]  ( .D(n325), .CP(Clk_s), .SD(Rst_n), .Q(n324) );
  FD4QM1P \receivedPacket_reg[19]  ( .D(n327), .CP(Clk_s), .SD(Rst_n), .Q(n326) );
  FD4QM1P \receivedPacket_reg[20]  ( .D(n329), .CP(Clk_s), .SD(Rst_n), .Q(n328) );
  FD4QM1P \receivedPacket_reg[21]  ( .D(n331), .CP(Clk_s), .SD(Rst_n), .Q(n330) );
  FD4QM1P \receivedPacket_reg[22]  ( .D(n333), .CP(Clk_s), .SD(Rst_n), .Q(n332) );
  FD4QM1P \receivedPacket_reg[23]  ( .D(n335), .CP(Clk_s), .SD(Rst_n), .Q(n334) );
  FD4QM1P \receivedPacket_reg[24]  ( .D(n337), .CP(Clk_s), .SD(Rst_n), .Q(n336) );
  FD4QM1P \receivedPacket_reg[25]  ( .D(n339), .CP(Clk_s), .SD(Rst_n), .Q(n338) );
  FD4QM1P \receivedPacket_reg[26]  ( .D(n341), .CP(Clk_s), .SD(Rst_n), .Q(n340) );
  FD4QM1P \receivedPacket_reg[27]  ( .D(n343), .CP(Clk_s), .SD(Rst_n), .Q(n342) );
  FD4QM1P \receivedPacket_reg[29]  ( .D(n347), .CP(Clk_s), .SD(Rst_n), .Q(n346) );
  FD4QM1P \receivedPacket_reg[31]  ( .D(n351), .CP(Clk_s), .SD(Rst_n), .Q(n350) );
  FD4QM1P \receivedPacket_reg[32]  ( .D(n353), .CP(Clk_s), .SD(Rst_n), .Q(n352) );
  FD2QM1P \RxData_reg[28]  ( .D(n277), .CP(Clk_s), .CD(Rst_n), .Q(RxData[28])
         );
  FD2QM1P \RxData_reg[17]  ( .D(n266), .CP(Clk_s), .CD(Rst_n), .Q(RxData[17])
         );
  FD4QM1P \receivedPacket_reg[28]  ( .D(n345), .CP(Clk_s), .SD(Rst_n), .Q(n344) );
  FD4QM1P \receivedPacket_reg[30]  ( .D(n349), .CP(Clk_s), .SD(Rst_n), .Q(n348) );
  FD2QM3P \RxData_reg[7]  ( .D(n256), .CP(Clk_s), .CD(Rst_n), .Q(RxData[7]) );
  FD2QM3P \RxData_reg[11]  ( .D(n260), .CP(Clk_s), .CD(Rst_n), .Q(RxData[11])
         );
  FD2QM3P \RxData_reg[18]  ( .D(n267), .CP(Clk_s), .CD(Rst_n), .Q(RxData[18])
         );
  FD2QM3P \RxData_reg[25]  ( .D(n274), .CP(Clk_s), .CD(Rst_n), .Q(RxData[25])
         );
  FD2QM3P \RxData_reg[30]  ( .D(n279), .CP(Clk_s), .CD(Rst_n), .Q(RxData[30])
         );
  FD2QM3P \RxData_reg[2]  ( .D(n251), .CP(Clk_s), .CD(Rst_n), .Q(RxData[2]) );
  FD2QM3P \RxData_reg[5]  ( .D(n254), .CP(Clk_s), .CD(Rst_n), .Q(RxData[5]) );
  FD2QM3P \RxData_reg[6]  ( .D(n255), .CP(Clk_s), .CD(Rst_n), .Q(RxData[6]) );
  FD2QM3P \RxData_reg[9]  ( .D(n258), .CP(Clk_s), .CD(Rst_n), .Q(RxData[9]) );
  FD2QM3P \RxData_reg[12]  ( .D(n261), .CP(Clk_s), .CD(Rst_n), .Q(RxData[12])
         );
  FD2QM3P \RxData_reg[15]  ( .D(n264), .CP(Clk_s), .CD(Rst_n), .Q(RxData[15])
         );
  FD2QM3P \RxData_reg[20]  ( .D(n269), .CP(Clk_s), .CD(Rst_n), .Q(RxData[20])
         );
  FD2QM3P \RxData_reg[23]  ( .D(n272), .CP(Clk_s), .CD(Rst_n), .Q(RxData[23])
         );
  FD2QM3P \RxData_reg[0]  ( .D(n249), .CP(Clk_s), .CD(Rst_n), .Q(RxData[0]) );
  FD2QM3P \RxData_reg[1]  ( .D(n250), .CP(Clk_s), .CD(Rst_n), .Q(RxData[1]) );
  FD2QM3P \RxData_reg[3]  ( .D(n252), .CP(Clk_s), .CD(Rst_n), .Q(RxData[3]) );
  FD2QM3P \RxData_reg[4]  ( .D(n253), .CP(Clk_s), .CD(Rst_n), .Q(RxData[4]) );
  FD2QM3P \RxData_reg[8]  ( .D(n257), .CP(Clk_s), .CD(Rst_n), .Q(RxData[8]) );
  FD2QM3P \RxData_reg[10]  ( .D(n259), .CP(Clk_s), .CD(Rst_n), .Q(RxData[10])
         );
  FD2QM3P \RxData_reg[13]  ( .D(n262), .CP(Clk_s), .CD(Rst_n), .Q(RxData[13])
         );
  FD2QM3P \RxData_reg[14]  ( .D(n263), .CP(Clk_s), .CD(Rst_n), .Q(RxData[14])
         );
  FD2QM3P \RxData_reg[16]  ( .D(n265), .CP(Clk_s), .CD(Rst_n), .Q(RxData[16])
         );
  FD2QM3P \RxData_reg[19]  ( .D(n268), .CP(Clk_s), .CD(Rst_n), .Q(RxData[19])
         );
  FD2QM3P \RxData_reg[21]  ( .D(n270), .CP(Clk_s), .CD(Rst_n), .Q(RxData[21])
         );
  FD2QM3P \RxData_reg[22]  ( .D(n271), .CP(Clk_s), .CD(Rst_n), .Q(RxData[22])
         );
  FD2QM3P \RxData_reg[24]  ( .D(n273), .CP(Clk_s), .CD(Rst_n), .Q(RxData[24])
         );
  FD2QM3P \RxData_reg[27]  ( .D(n276), .CP(Clk_s), .CD(Rst_n), .Q(RxData[27])
         );
  FD2QM3P \RxData_reg[29]  ( .D(n278), .CP(Clk_s), .CD(Rst_n), .Q(RxData[29])
         );
  FD2QM3P \RxData_reg[31]  ( .D(n280), .CP(Clk_s), .CD(Rst_n), .Q(RxData[31])
         );
  FD2QM3P \RxData_reg[26]  ( .D(n275), .CP(Clk_s), .CD(Rst_n), .Q(RxData[26])
         );
  FD2QM1P \zeroCounter_reg[0]  ( .D(N24), .CP(Clk_s), .CD(Rst_n), .Q(
        zeroCounter[0]) );
  FD2QM1P Rx_Ready_reg ( .D(N27), .CP(Clk_s), .CD(Rst_n), .Q(Rx_Ready) );
  FD2QM1P \zeroCounter_reg[1]  ( .D(N25), .CP(Clk_s), .CD(Rst_n), .Q(
        zeroCounter[1]) );
  FD2QM1P \zeroCounter_reg[2]  ( .D(N26), .CP(Clk_s), .CD(Rst_n), .Q(
        zeroCounter[2]) );
  FD2QM1P bitStuff_reg ( .D(N22), .CP(Clk_s), .CD(Rst_n), .Q(bitStuff) );
  FD2QM1P dataRx_reg ( .D(n247), .CP(Clk_s), .CD(Rst_n), .Q(dataRx) );
  FD2QM1P \receivedCounter_reg[0]  ( .D(n248), .CP(Clk_s), .CD(Rst_n), .Q(
        receivedCounter[0]) );
  FD2QM1P Rx_Error_reg ( .D(N229), .CP(Clk_s), .CD(Rst_n), .Q(Rx_Error) );
  FD2QM1P bufferFull_reg ( .D(N242), .CP(Clk_s), .CD(Rst_n), .Q(bufferFull) );
  FD2QM1P \receivedCounter_reg[1]  ( .D(n281), .CP(Clk_s), .CD(Rst_n), .Q(
        receivedCounter[1]) );
  FD2QM1P \receivedCounter_reg[3]  ( .D(n283), .CP(Clk_s), .CD(Rst_n), .Q(
        receivedCounter[3]) );
  FD2QM1P \receivedCounter_reg[2]  ( .D(n282), .CP(Clk_s), .CD(Rst_n), .Q(
        receivedCounter[2]) );
  FD2QM1P RxData_Valid_reg ( .D(N243), .CP(Clk_s), .CD(Rst_n), .Q(RxData_Valid) );
  FD2QM1P \receivedCounter_reg[4]  ( .D(n284), .CP(Clk_s), .CD(Rst_n), .Q(
        receivedCounter[4]) );
  FD2QM1P \receivedCounter_reg[5]  ( .D(n285), .CP(Clk_s), .CD(Rst_n), .Q(
        receivedCounter[5]) );
  ND2M1P U3 ( .A(n117), .B(n115), .Z(n79) );
  N1M3P U4 ( .A(n79), .Z(n80) );
  N1M4P U5 ( .A(n81), .Z(n75) );
  MUX21LM1P U6 ( .A(n324), .B(n135), .S(n78), .Z(n266) );
  ENFM1P U7 ( .A(n310), .B(n308), .Z(n74) );
  EN3M1P U8 ( .A(n312), .B(n298), .C(n74), .Z(n103) );
  AOI22DNM1P U9 ( .A(n152), .B(n80), .D(n352), .C(n75), .Z(n353) );
  N1M12P U10 ( .A(n77), .Z(n76) );
  NR2FM2P U11 ( .A(n116), .B(n115), .Z(n206) );
  OAI21M2P U12 ( .A(n84), .B(n83), .C(receivedCounter[5]), .Z(n115) );
  ND2M1P U13 ( .A(dataRx), .B(n286), .Z(n225) );
  N1M1P U14 ( .A(bufferFull), .Z(n227) );
  N1M2P U15 ( .A(n344), .Z(n243) );
  N1M6P U16 ( .A(n149), .Z(n77) );
  N1M6P U17 ( .A(n77), .Z(n78) );
  ND2FM3P U18 ( .A(n206), .B(n117), .Z(n149) );
  MUX21LFM1P U19 ( .A(n346), .B(n146), .S(n76), .Z(n277) );
  ND2FM2P U20 ( .A(n113), .B(n227), .Z(n116) );
  NR2FM1P U21 ( .A(n225), .B(bitStuff), .Z(n117) );
  N1M1P U22 ( .A(n348), .Z(n245) );
  N1M1P U23 ( .A(n342), .Z(n242) );
  OR2M1P U24 ( .A(receivedCounter[3]), .B(receivedCounter[0]), .Z(n83) );
  NR2BNM1P U25 ( .B(n117), .A(n115), .Z(n114) );
  ND2BNM1P U26 ( .B(receivedCounter[1]), .A(n82), .Z(n84) );
  AND3M1P U27 ( .A(n116), .B(n114), .C(n227), .Z(N229) );
  AOI22M1P U28 ( .A(n152), .B(n75), .C(n245), .D(n80), .Z(n351) );
  N1M1P U29 ( .A(n332), .Z(n209) );
  N1M1P U30 ( .A(n340), .Z(n213) );
  N1M1P U31 ( .A(n334), .Z(n210) );
  N1M1P U32 ( .A(n338), .Z(n212) );
  N1M1P U33 ( .A(n336), .Z(n211) );
  AOI22M1P U34 ( .A(n208), .B(n75), .C(n80), .D(n153), .Z(n331) );
  N1M1P U35 ( .A(n330), .Z(n208) );
  OAI21M1P U36 ( .A(n227), .B(n220), .C(n207), .Z(N242) );
  N1M1P U37 ( .A(n206), .Z(n207) );
  NR2BNM1P U38 ( .B(RxData_Valid), .A(n206), .Z(n151) );
  N1M1P U39 ( .A(receivedCounter[3]), .Z(n216) );
  AOI22M1P U40 ( .A(n205), .B(n75), .C(n241), .D(S_Data), .Z(n289) );
  AOI22M1P U41 ( .A(n157), .B(n75), .C(n80), .D(n190), .Z(n321) );
  AOI22M1P U42 ( .A(n204), .B(n75), .C(n80), .D(n205), .Z(n291) );
  N1M1P U43 ( .A(n288), .Z(n205) );
  AOI22M1P U44 ( .A(n203), .B(n75), .C(n80), .D(n204), .Z(n293) );
  N1M1P U45 ( .A(n290), .Z(n204) );
  AOI22M1P U46 ( .A(n202), .B(n75), .C(n80), .D(n203), .Z(n295) );
  N1M1P U47 ( .A(n292), .Z(n203) );
  AOI22M1P U48 ( .A(n194), .B(n75), .C(n80), .D(n195), .Z(n311) );
  AOI22M1P U49 ( .A(n155), .B(n75), .C(n80), .D(n156), .Z(n325) );
  AOI22M1P U50 ( .A(n191), .B(n75), .C(n80), .D(n192), .Z(n317) );
  AOI22M1P U51 ( .A(n193), .B(n75), .C(n80), .D(n194), .Z(n313) );
  N1M1P U52 ( .A(n310), .Z(n194) );
  AOI22M1P U53 ( .A(n195), .B(n75), .C(n80), .D(n196), .Z(n309) );
  N1M1P U54 ( .A(n308), .Z(n195) );
  AOI22M1P U55 ( .A(n153), .B(n75), .C(n80), .D(n154), .Z(n329) );
  N1M1P U56 ( .A(n328), .Z(n153) );
  N1M1P U57 ( .A(n350), .Z(n152) );
  AOI22M1P U58 ( .A(n196), .B(n75), .C(n80), .D(n197), .Z(n307) );
  N1M1P U59 ( .A(n306), .Z(n196) );
  AOI22M1P U60 ( .A(n198), .B(n75), .C(n80), .D(n199), .Z(n303) );
  AOI22M1P U61 ( .A(n154), .B(n75), .C(n80), .D(n155), .Z(n327) );
  N1M1P U62 ( .A(n326), .Z(n154) );
  AOI22M1P U63 ( .A(n192), .B(n75), .C(n80), .D(n193), .Z(n315) );
  N1M1P U64 ( .A(n312), .Z(n193) );
  N1M1P U65 ( .A(n314), .Z(n192) );
  AOI22M1P U66 ( .A(n201), .B(n75), .C(n80), .D(n202), .Z(n297) );
  N1M1P U67 ( .A(n294), .Z(n202) );
  AOI22M1P U68 ( .A(n199), .B(n75), .C(n80), .D(n200), .Z(n301) );
  N1M1P U69 ( .A(n300), .Z(n199) );
  AOI22M1P U70 ( .A(n200), .B(n75), .C(n80), .D(n201), .Z(n299) );
  N1M1P U71 ( .A(n296), .Z(n201) );
  N1M1P U72 ( .A(n298), .Z(n200) );
  AOI22M1P U73 ( .A(n156), .B(n75), .C(n80), .D(n157), .Z(n323) );
  N1M1P U74 ( .A(n320), .Z(n157) );
  N1M1P U75 ( .A(n322), .Z(n156) );
  AOI22M1P U76 ( .A(n197), .B(n75), .C(n80), .D(n198), .Z(n305) );
  N1M1P U77 ( .A(n302), .Z(n198) );
  N1M1P U78 ( .A(n304), .Z(n197) );
  AOI22M1P U79 ( .A(n190), .B(n75), .C(n80), .D(n191), .Z(n319) );
  N1M1P U80 ( .A(n316), .Z(n191) );
  N1M1P U81 ( .A(n318), .Z(n190) );
  N1M1P U82 ( .A(receivedCounter[4]), .Z(n215) );
  ND2BNM1P U83 ( .B(n227), .A(n114), .Z(n85) );
  N1M1P U84 ( .A(receivedCounter[0]), .Z(n214) );
  N1M1P U85 ( .A(receivedCounter[2]), .Z(n217) );
  N1M1P U86 ( .A(RxData[17]), .Z(n135) );
  MUX21LM1P U87 ( .A(n344), .B(n145), .S(n78), .Z(n276) );
  N1M1P U88 ( .A(RxData[27]), .Z(n145) );
  MUX21LM1P U89 ( .A(n290), .B(n118), .S(n76), .Z(n249) );
  N1M1P U90 ( .A(RxData[0]), .Z(n118) );
  MUX21LM1P U91 ( .A(n310), .B(n128), .S(n78), .Z(n259) );
  N1M1P U92 ( .A(RxData[10]), .Z(n128) );
  MUX21LM1P U93 ( .A(n306), .B(n126), .S(n76), .Z(n257) );
  N1M1P U94 ( .A(RxData[8]), .Z(n126) );
  MUX21LM1P U95 ( .A(n328), .B(n137), .S(n76), .Z(n268) );
  N1M1P U96 ( .A(RxData[19]), .Z(n137) );
  MUX21LM1P U97 ( .A(n334), .B(n140), .S(n78), .Z(n271) );
  N1M1P U98 ( .A(RxData[22]), .Z(n140) );
  MUX21LM1P U99 ( .A(n332), .B(n139), .S(n76), .Z(n270) );
  N1M1P U100 ( .A(RxData[21]), .Z(n139) );
  MUX21LM1P U101 ( .A(n338), .B(n142), .S(n76), .Z(n273) );
  N1M1P U102 ( .A(RxData[24]), .Z(n142) );
  MUX21LM1P U103 ( .A(n352), .B(n150), .S(n78), .Z(n280) );
  N1M1P U104 ( .A(RxData[31]), .Z(n150) );
  MUX21LM1P U105 ( .A(n316), .B(n131), .S(n76), .Z(n262) );
  N1M1P U106 ( .A(RxData[13]), .Z(n131) );
  MUX21LM1P U107 ( .A(n322), .B(n134), .S(n76), .Z(n265) );
  N1M1P U108 ( .A(RxData[16]), .Z(n134) );
  MUX21LM1P U109 ( .A(n296), .B(n121), .S(n76), .Z(n252) );
  N1M1P U110 ( .A(RxData[3]), .Z(n121) );
  MUX21LM1P U111 ( .A(n298), .B(n122), .S(n76), .Z(n253) );
  N1M1P U112 ( .A(RxData[4]), .Z(n122) );
  MUX21LM1P U113 ( .A(n292), .B(n119), .S(n78), .Z(n250) );
  N1M1P U114 ( .A(RxData[1]), .Z(n119) );
  MUX21LM1P U115 ( .A(n318), .B(n132), .S(n76), .Z(n263) );
  N1M1P U116 ( .A(RxData[14]), .Z(n132) );
  MUX21LM1P U117 ( .A(n342), .B(n144), .S(n76), .Z(n275) );
  N1M1P U118 ( .A(RxData[26]), .Z(n144) );
  MUX21LM1P U119 ( .A(n300), .B(n123), .S(n78), .Z(n254) );
  N1M1P U120 ( .A(RxData[5]), .Z(n123) );
  MUX21LM1P U121 ( .A(n302), .B(n124), .S(n76), .Z(n255) );
  N1M1P U122 ( .A(RxData[6]), .Z(n124) );
  MUX21LM1P U123 ( .A(n336), .B(n141), .S(n76), .Z(n272) );
  N1M1P U124 ( .A(RxData[23]), .Z(n141) );
  MUX21LM1P U125 ( .A(n308), .B(n127), .S(n78), .Z(n258) );
  N1M1P U126 ( .A(RxData[9]), .Z(n127) );
  MUX21LM1P U127 ( .A(n294), .B(n120), .S(n76), .Z(n251) );
  N1M1P U128 ( .A(RxData[2]), .Z(n120) );
  MUX21LM1P U129 ( .A(n330), .B(n138), .S(n78), .Z(n269) );
  N1M1P U130 ( .A(RxData[20]), .Z(n138) );
  MUX21LM1P U131 ( .A(n314), .B(n130), .S(n76), .Z(n261) );
  N1M1P U132 ( .A(RxData[12]), .Z(n130) );
  MUX21LM1P U133 ( .A(n320), .B(n133), .S(n78), .Z(n264) );
  N1M1P U134 ( .A(RxData[15]), .Z(n133) );
  MUX21LM1P U135 ( .A(n326), .B(n136), .S(n76), .Z(n267) );
  N1M1P U136 ( .A(RxData[18]), .Z(n136) );
  MUX21LM1P U137 ( .A(n350), .B(n148), .S(n78), .Z(n279) );
  N1M1P U138 ( .A(RxData[30]), .Z(n148) );
  MUX21LM1P U139 ( .A(n304), .B(n125), .S(n76), .Z(n256) );
  N1M1P U140 ( .A(RxData[7]), .Z(n125) );
  MUX21LM1P U141 ( .A(n340), .B(n143), .S(n76), .Z(n274) );
  N1M1P U142 ( .A(RxData[25]), .Z(n143) );
  MUX21LM1P U143 ( .A(n312), .B(n129), .S(n76), .Z(n260) );
  N1M1P U144 ( .A(RxData[11]), .Z(n129) );
  N1M1P U145 ( .A(RxData[28]), .Z(n146) );
  MUX21LM1P U146 ( .A(n348), .B(n147), .S(n76), .Z(n278) );
  NR2M1P U147 ( .A(receivedCounter[2]), .B(receivedCounter[4]), .Z(n82) );
  ENFM1P U148 ( .A(n112), .B(n111), .Z(n113) );
  ENFM1P U149 ( .A(n110), .B(n109), .Z(n111) );
  EOFM1P U150 ( .A(n108), .B(n107), .Z(n109) );
  EOFM1P U151 ( .A(n219), .B(n106), .Z(n107) );
  ENFM1P U152 ( .A(n155), .B(n105), .Z(n106) );
  ENFM1P U153 ( .A(n332), .B(n336), .Z(n105) );
  N1M1P U154 ( .A(n324), .Z(n155) );
  AOI22M1P U155 ( .A(n348), .B(n346), .C(n244), .D(n245), .Z(n219) );
  N1M1P U156 ( .A(n346), .Z(n244) );
  EOFM1P U157 ( .A(n104), .B(n218), .Z(n108) );
  AOI22M1P U158 ( .A(n344), .B(n342), .C(n242), .D(n243), .Z(n218) );
  EOFM1P U159 ( .A(n328), .B(n326), .Z(n104) );
  ENFM1P U160 ( .A(n103), .B(n102), .Z(n110) );
  ENFM1P U161 ( .A(n101), .B(n100), .Z(n102) );
  ENFM1P U162 ( .A(n322), .B(n320), .Z(n100) );
  ENFM1P U163 ( .A(n318), .B(n300), .Z(n101) );
  ENFM1P U164 ( .A(n99), .B(n98), .Z(n112) );
  ENFM1P U165 ( .A(n97), .B(n96), .Z(n98) );
  ENFM1P U166 ( .A(n95), .B(n94), .Z(n96) );
  EOFM1P U167 ( .A(n306), .B(n304), .Z(n94) );
  ENFM1P U168 ( .A(n296), .B(n302), .Z(n95) );
  ENFM1P U169 ( .A(n93), .B(n92), .Z(n97) );
  EOFM1P U170 ( .A(n292), .B(n350), .Z(n92) );
  ENFM1P U171 ( .A(n290), .B(n294), .Z(n93) );
  ENFM1P U172 ( .A(n91), .B(n90), .Z(n99) );
  ENFM1P U173 ( .A(n89), .B(n88), .Z(n90) );
  ENFM1P U174 ( .A(n316), .B(n314), .Z(n88) );
  ENFM1P U175 ( .A(n352), .B(n288), .Z(n89) );
  ENFM1P U176 ( .A(n87), .B(n86), .Z(n91) );
  ENFM1P U177 ( .A(n338), .B(n330), .Z(n86) );
  EOFM1P U178 ( .A(n334), .B(n340), .Z(n87) );
  N1M1P U179 ( .A(RxData[29]), .Z(n147) );
  N1M2P U180 ( .A(n246), .Z(n81) );
  OAI21M1P U181 ( .A(n225), .B(n226), .C(n85), .Z(n246) );
  OA21M1P U182 ( .A(n151), .B(bufferFull), .C(Core_Rcv_Ready), .Z(N243) );
  ND2M1P U183 ( .A(zeroCounter[1]), .B(zeroCounter[0]), .Z(n221) );
  NR3M1P U184 ( .A(S_Data), .B(zeroCounter[2]), .C(n221), .Z(N26) );
  N1M1P U185 ( .A(receivedCounter[5]), .Z(n239) );
  AND2M1P U186 ( .A(N26), .B(n239), .Z(N22) );
  NR3M1P U187 ( .A(S_Data), .B(zeroCounter[2]), .C(zeroCounter[0]), .Z(N24) );
  NR2BNM1P U188 ( .B(RxData_Valid), .A(Core_Rcv_Ready), .Z(n220) );
  OAI21M1P U189 ( .A(zeroCounter[1]), .B(zeroCounter[0]), .C(n221), .Z(n222)
         );
  NR3M1P U190 ( .A(S_Data), .B(zeroCounter[2]), .C(n222), .Z(N25) );
  NR2BNM1P U191 ( .B(n286), .A(dataRx), .Z(N27) );
  ND2M1P U192 ( .A(n286), .B(n79), .Z(n241) );
  N1M1P U193 ( .A(bitStuff), .Z(n226) );
  ND2BNM1P U194 ( .B(n241), .A(n81), .Z(n247) );
  ND2M1P U195 ( .A(n80), .B(n214), .Z(n228) );
  OAI211M1P U196 ( .A(n81), .B(n214), .C(n286), .D(n228), .Z(n248) );
  AOI21M1P U197 ( .A(n80), .B(n214), .C(n75), .Z(n229) );
  N1M1P U198 ( .A(receivedCounter[1]), .Z(n233) );
  NR2M1P U199 ( .A(receivedCounter[1]), .B(n79), .Z(n230) );
  OAI22CDNM1P U200 ( .A(n229), .B(n233), .C(receivedCounter[0]), .D(n230), .Z(
        n281) );
  AOI211M1P U201 ( .A(n80), .B(n214), .C(n230), .D(n75), .Z(n232) );
  ND3M1P U202 ( .A(receivedCounter[1]), .B(receivedCounter[0]), .C(n80), .Z(
        n231) );
  AOI22M1P U203 ( .A(receivedCounter[2]), .B(n232), .C(n231), .D(n217), .Z(
        n282) );
  NR3M1P U204 ( .A(n233), .B(n217), .C(n214), .Z(n237) );
  N1M1P U205 ( .A(n237), .Z(n234) );
  AOI21M1P U206 ( .A(n234), .B(n80), .C(n75), .Z(n236) );
  ND2M1P U207 ( .A(n80), .B(n216), .Z(n235) );
  OAI22M1P U208 ( .A(n236), .B(n216), .C(n235), .D(n234), .Z(n283) );
  OA21M1P U209 ( .A(n79), .B(receivedCounter[3]), .C(n236), .Z(n240) );
  ND3M1P U210 ( .A(receivedCounter[3]), .B(n80), .C(n237), .Z(n238) );
  AOI22M1P U211 ( .A(receivedCounter[4]), .B(n240), .C(n238), .D(n215), .Z(
        n284) );
  OAI22M1P U212 ( .A(n240), .B(n239), .C(n215), .D(n238), .Z(n285) );
  ND2BNM1P U213 ( .B(S_Data), .A(zeroCounter[2]), .Z(n287) );
  AOI22M1P U214 ( .A(n80), .B(n208), .C(n209), .D(n75), .Z(n333) );
  AOI22M1P U215 ( .A(n80), .B(n209), .C(n210), .D(n75), .Z(n335) );
  AOI22M1P U216 ( .A(n80), .B(n210), .C(n211), .D(n75), .Z(n337) );
  AOI22M1P U217 ( .A(n80), .B(n211), .C(n212), .D(n75), .Z(n339) );
  AOI22M1P U218 ( .A(n80), .B(n212), .C(n213), .D(n75), .Z(n341) );
  AOI22M1P U219 ( .A(n80), .B(n213), .C(n242), .D(n75), .Z(n343) );
  AOI22M1P U220 ( .A(n80), .B(n242), .C(n243), .D(n75), .Z(n345) );
  AOI22M1P U221 ( .A(n80), .B(n243), .C(n244), .D(n75), .Z(n347) );
  AOI22M1P U222 ( .A(n80), .B(n244), .C(n245), .D(n75), .Z(n349) );
endmodule


module tx_1 ( Clk_s, Rst_n, TxData_Valid, TxData, Error_Ack, Rx_Ready, 
        Rx_Error, Tx_Ready, Tx_Error, S_Data );
  input [31:0] TxData;
  input Clk_s, Rst_n, TxData_Valid, Error_Ack, Rx_Ready, Rx_Error;
  output Tx_Ready, Tx_Error, S_Data;
  wire   N100, N101, N102, N103, N104, N105, N106, N107, N108, N109, N110,
         N111, N112, N113, N114, N115, N116, N117, N118, N119, N120, N121,
         N122, N123, N124, N125, N126, N127, N128, N129, N130, N131, N132,
         N146, n17, n18, n19, n20, n21, n22, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167;
  wire   [32:0] transmissionPacket;
  wire   [5:0] bitCount;

  FD4QM1P zeroPatternDetected_reg ( .D(n154), .CP(Clk_s), .SD(Rst_n), .Q(n153)
         );
  FD4QM1P DataTxInProg_reg ( .D(n156), .CP(Clk_s), .SD(Rst_n), .Q(n155) );
  FD4QM1P Tx_Ready_reg ( .D(n143), .CP(Clk_s), .SD(Rst_n), .Q(Tx_Ready) );
  FD2LQM1P \transmissionPacket_reg[1]  ( .D(TxData[0]), .LD(n58), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[1]) );
  FD2LQM1P \transmissionPacket_reg[2]  ( .D(TxData[1]), .LD(n58), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[2]) );
  FD2LQM1P \transmissionPacket_reg[3]  ( .D(TxData[2]), .LD(n58), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[3]) );
  FD2LQM1P \transmissionPacket_reg[4]  ( .D(TxData[3]), .LD(n58), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[4]) );
  FD2LQM1P \transmissionPacket_reg[5]  ( .D(TxData[4]), .LD(n58), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[5]) );
  FD2LQM1P \transmissionPacket_reg[6]  ( .D(TxData[5]), .LD(n58), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[6]) );
  FD2LQM1P \transmissionPacket_reg[7]  ( .D(TxData[6]), .LD(n58), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[7]) );
  FD2LQM1P \transmissionPacket_reg[8]  ( .D(TxData[7]), .LD(n58), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[8]) );
  FD2LQM1P \transmissionPacket_reg[9]  ( .D(TxData[8]), .LD(n58), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[9]) );
  FD2LQM1P \transmissionPacket_reg[10]  ( .D(TxData[9]), .LD(n58), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[10]) );
  FD2LQM1P \transmissionPacket_reg[11]  ( .D(TxData[10]), .LD(n58), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[11]) );
  FD2LQM1P \transmissionPacket_reg[12]  ( .D(TxData[11]), .LD(n58), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[12]) );
  FD2LQM1P \transmissionPacket_reg[13]  ( .D(TxData[12]), .LD(n58), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[13]) );
  FD2LQM1P \transmissionPacket_reg[14]  ( .D(TxData[13]), .LD(n58), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[14]) );
  FD2LQM1P \transmissionPacket_reg[15]  ( .D(TxData[14]), .LD(n58), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[15]) );
  FD2LQM1P \transmissionPacket_reg[16]  ( .D(TxData[15]), .LD(n58), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[16]) );
  FD2LQM1P \transmissionPacket_reg[17]  ( .D(TxData[16]), .LD(n58), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[17]) );
  FD2LQM1P \transmissionPacket_reg[18]  ( .D(TxData[17]), .LD(n58), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[18]) );
  FD2LQM1P \transmissionPacket_reg[19]  ( .D(TxData[18]), .LD(n58), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[19]) );
  FD2LQM1P \transmissionPacket_reg[20]  ( .D(TxData[19]), .LD(n58), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[20]) );
  FD2LQM1P \transmissionPacket_reg[21]  ( .D(TxData[20]), .LD(n58), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[21]) );
  FD2LQM1P \transmissionPacket_reg[22]  ( .D(TxData[21]), .LD(n58), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[22]) );
  FD2LQM1P \transmissionPacket_reg[23]  ( .D(TxData[22]), .LD(n152), .CP(Clk_s), .CD(Rst_n), .Q(transmissionPacket[23]) );
  FD2LQM1P \transmissionPacket_reg[24]  ( .D(TxData[23]), .LD(n152), .CP(Clk_s), .CD(Rst_n), .Q(transmissionPacket[24]) );
  FD2LQM1P \transmissionPacket_reg[25]  ( .D(TxData[24]), .LD(n152), .CP(Clk_s), .CD(Rst_n), .Q(transmissionPacket[25]) );
  FD2LQM1P \transmissionPacket_reg[26]  ( .D(TxData[25]), .LD(n152), .CP(Clk_s), .CD(Rst_n), .Q(transmissionPacket[26]) );
  FD2LQM1P \transmissionPacket_reg[27]  ( .D(TxData[26]), .LD(n152), .CP(Clk_s), .CD(Rst_n), .Q(transmissionPacket[27]) );
  FD2LQM1P \transmissionPacket_reg[28]  ( .D(TxData[27]), .LD(n152), .CP(Clk_s), .CD(Rst_n), .Q(transmissionPacket[28]) );
  FD2LQM1P \transmissionPacket_reg[29]  ( .D(TxData[28]), .LD(n152), .CP(Clk_s), .CD(Rst_n), .Q(transmissionPacket[29]) );
  FD2LQM1P \transmissionPacket_reg[30]  ( .D(TxData[29]), .LD(n152), .CP(Clk_s), .CD(Rst_n), .Q(transmissionPacket[30]) );
  FD2LQM1P \transmissionPacket_reg[31]  ( .D(TxData[30]), .LD(n152), .CP(Clk_s), .CD(Rst_n), .Q(transmissionPacket[31]) );
  FD2LQM1P \transmissionPacket_reg[32]  ( .D(TxData[31]), .LD(n58), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[32]) );
  FD4QM1P \startSequenceCount_reg[1]  ( .D(n158), .CP(Clk_s), .SD(Rst_n), .Q(
        n157) );
  FD4QM1P \startSequenceCount_reg[2]  ( .D(n160), .CP(Clk_s), .SD(Rst_n), .Q(
        n159) );
  FD4QM1P \startSequenceCount_reg[0]  ( .D(n162), .CP(Clk_s), .SD(Rst_n), .Q(
        n161) );
  FD4QM1P startSequence_reg ( .D(n145), .CP(Clk_s), .SD(Rst_n), .Q(n163) );
  FD4QM1P \zeroCount_reg[0]  ( .D(n165), .CP(Clk_s), .SD(Rst_n), .Q(n164) );
  FD4QM1P \zeroCount_reg[1]  ( .D(n167), .CP(Clk_s), .SD(Rst_n), .Q(n166) );
  FD4QM1P S_Data_reg ( .D(N146), .CP(Clk_s), .SD(Rst_n), .Q(S_Data) );
  FD2QM1P \bitCount_reg[0]  ( .D(n151), .CP(Clk_s), .CD(Rst_n), .Q(bitCount[0]) );
  FD2QM1P \bitCount_reg[3]  ( .D(n148), .CP(Clk_s), .CD(Rst_n), .Q(bitCount[3]) );
  FD2QM1P \bitCount_reg[1]  ( .D(n150), .CP(Clk_s), .CD(Rst_n), .Q(bitCount[1]) );
  FD2QM1P \bitCount_reg[4]  ( .D(n147), .CP(Clk_s), .CD(Rst_n), .Q(bitCount[4]) );
  FD2QM1P \bitCount_reg[5]  ( .D(n146), .CP(Clk_s), .CD(Rst_n), .Q(bitCount[5]) );
  FD2QM1P \bitCount_reg[2]  ( .D(n149), .CP(Clk_s), .CD(Rst_n), .Q(bitCount[2]) );
  FD2QM1P \transmissionPacket_reg[0]  ( .D(n144), .CP(Clk_s), .CD(Rst_n), .Q(
        transmissionPacket[0]) );
  NR2BNM1P U3 ( .B(bitCount[4]), .A(bitCount[5]), .Z(n46) );
  ND2M1P U4 ( .A(bitCount[1]), .B(bitCount[0]), .Z(n53) );
  ND2BNM1P U5 ( .B(bitCount[1]), .A(bitCount[0]), .Z(n55) );
  OR2M1P U6 ( .A(bitCount[0]), .B(bitCount[1]), .Z(n54) );
  N1M1P U7 ( .A(bitCount[2]), .Z(n124) );
  ND4M1P U8 ( .A(n153), .B(n163), .C(n138), .D(n81), .Z(n131) );
  AND2M1P U9 ( .A(Tx_Ready), .B(TxData_Valid), .Z(n152) );
  AOI22DNM1P U10 ( .A(n166), .B(n142), .D(n140), .C(n141), .Z(n17) );
  OA21M1P U11 ( .A(n166), .B(n20), .C(n17), .Z(n167) );
  N1M1P U12 ( .A(n131), .Z(n133) );
  NR3M1P U13 ( .A(n37), .B(n36), .C(n35), .Z(n40) );
  ND2BNM2P U14 ( .B(bitCount[0]), .A(bitCount[1]), .Z(n18) );
  BUFM2P U15 ( .A(n152), .Z(n58) );
  ND2BNM1P U16 ( .B(n19), .A(n164), .Z(n20) );
  NR2M1P U17 ( .A(n19), .B(n164), .Z(n142) );
  N1M1P U18 ( .A(bitCount[3]), .Z(n57) );
  ND2M1P U19 ( .A(n48), .B(n46), .Z(n43) );
  OA21M1P U20 ( .A(n164), .B(n140), .C(n20), .Z(n165) );
  NR2M1P U21 ( .A(n18), .B(n52), .Z(N106) );
  NR2M1P U22 ( .A(n18), .B(n47), .Z(N130) );
  NR2M1P U23 ( .A(n50), .B(n18), .Z(N102) );
  NR2M1P U24 ( .A(n18), .B(n45), .Z(N126) );
  NR2M1P U25 ( .A(n18), .B(n44), .Z(N122) );
  NR2M1P U26 ( .A(n18), .B(n43), .Z(N118) );
  NR2M1P U27 ( .A(n18), .B(n42), .Z(N114) );
  NR2M1P U28 ( .A(n56), .B(n18), .Z(N110) );
  ND2M1P U29 ( .A(n41), .B(n40), .Z(n19) );
  AOI22M1P U30 ( .A(transmissionPacket[13]), .B(N119), .C(
        transmissionPacket[12]), .D(N120), .Z(n21) );
  AOI22M1P U31 ( .A(transmissionPacket[22]), .B(N110), .C(
        transmissionPacket[21]), .D(N111), .Z(n22) );
  AOI22M1P U32 ( .A(transmissionPacket[23]), .B(N109), .C(
        transmissionPacket[20]), .D(N112), .Z(n29) );
  AOI22M1P U33 ( .A(transmissionPacket[2]), .B(N130), .C(transmissionPacket[1]), .D(N131), .Z(n30) );
  AOI22M1P U34 ( .A(transmissionPacket[4]), .B(N128), .C(transmissionPacket[6]), .D(N126), .Z(n31) );
  AOI22M1P U35 ( .A(transmissionPacket[5]), .B(N127), .C(transmissionPacket[3]), .D(N129), .Z(n32) );
  AOI22M1P U36 ( .A(transmissionPacket[7]), .B(N125), .C(transmissionPacket[9]), .D(N123), .Z(n33) );
  AOI22M1P U37 ( .A(transmissionPacket[11]), .B(N121), .C(
        transmissionPacket[10]), .D(N122), .Z(n34) );
  ND4M1P U38 ( .A(n69), .B(n68), .C(n67), .D(n21), .Z(n35) );
  ND4M1P U39 ( .A(n65), .B(n64), .C(n29), .D(n22), .Z(n36) );
  ND4M1P U40 ( .A(n30), .B(n60), .C(n59), .D(n66), .Z(n37) );
  ND4M1P U41 ( .A(n34), .B(n33), .C(n32), .D(n31), .Z(n38) );
  ND3M1P U42 ( .A(n138), .B(n153), .C(n163), .Z(n39) );
  AOI211M1P U43 ( .A(N124), .B(transmissionPacket[8]), .C(n39), .D(n38), .Z(
        n41) );
  NR2M1P U44 ( .A(n54), .B(n50), .Z(N100) );
  NR2M1P U45 ( .A(n56), .B(n53), .Z(N111) );
  NR2M1P U46 ( .A(n54), .B(n42), .Z(N112) );
  NR2M1P U47 ( .A(n42), .B(n55), .Z(N113) );
  NR2M1P U48 ( .A(n53), .B(n42), .Z(N115) );
  NR2M1P U49 ( .A(n54), .B(n43), .Z(N116) );
  NR2M1P U50 ( .A(n55), .B(n43), .Z(N117) );
  NR2M1P U51 ( .A(n53), .B(n43), .Z(N119) );
  NR2M1P U52 ( .A(n50), .B(n55), .Z(N101) );
  NR2M1P U53 ( .A(n54), .B(n44), .Z(N120) );
  NR2M1P U54 ( .A(n55), .B(n44), .Z(N121) );
  NR2M1P U55 ( .A(n53), .B(n44), .Z(N123) );
  NR2M1P U56 ( .A(n54), .B(n45), .Z(N124) );
  NR2M1P U57 ( .A(n55), .B(n45), .Z(N125) );
  NR2M1P U58 ( .A(n53), .B(n45), .Z(N127) );
  NR2M1P U59 ( .A(n54), .B(n47), .Z(N128) );
  NR2M1P U60 ( .A(n55), .B(n47), .Z(N129) );
  NR2M1P U61 ( .A(n53), .B(n47), .Z(N131) );
  NR3M1P U62 ( .A(bitCount[4]), .B(n54), .C(n49), .Z(N132) );
  NR2M1P U63 ( .A(n50), .B(n53), .Z(N103) );
  NR2M1P U64 ( .A(n54), .B(n52), .Z(N104) );
  NR2M1P U65 ( .A(n55), .B(n52), .Z(N105) );
  NR2M1P U66 ( .A(n53), .B(n52), .Z(N107) );
  NR2M1P U67 ( .A(n54), .B(n56), .Z(N108) );
  NR2M1P U68 ( .A(n56), .B(n55), .Z(N109) );
  NR2M1P U69 ( .A(bitCount[5]), .B(bitCount[4]), .Z(n51) );
  NR2M1P U70 ( .A(bitCount[2]), .B(bitCount[3]), .Z(n48) );
  ND2M1P U71 ( .A(n51), .B(n48), .Z(n50) );
  ND3M1P U72 ( .A(n51), .B(bitCount[3]), .C(n124), .Z(n56) );
  ND3M1P U73 ( .A(n51), .B(bitCount[2]), .C(bitCount[3]), .Z(n42) );
  ND3M1P U74 ( .A(bitCount[2]), .B(n46), .C(n57), .Z(n44) );
  ND3M1P U75 ( .A(bitCount[3]), .B(n46), .C(n124), .Z(n45) );
  ND3M1P U76 ( .A(bitCount[2]), .B(bitCount[3]), .C(n46), .Z(n47) );
  ND2M1P U77 ( .A(bitCount[5]), .B(n48), .Z(n49) );
  ND3M1P U78 ( .A(bitCount[2]), .B(n51), .C(n57), .Z(n52) );
  AOI22M1P U79 ( .A(transmissionPacket[5]), .B(N127), .C(transmissionPacket[3]), .D(N129), .Z(n62) );
  AOI22M1P U80 ( .A(transmissionPacket[2]), .B(N130), .C(transmissionPacket[1]), .D(N131), .Z(n61) );
  AOI22M1P U81 ( .A(transmissionPacket[32]), .B(N100), .C(
        transmissionPacket[0]), .D(N132), .Z(n60) );
  AOI22M1P U82 ( .A(transmissionPacket[30]), .B(N102), .C(
        transmissionPacket[31]), .D(N101), .Z(n59) );
  ND4M1P U83 ( .A(n62), .B(n61), .C(n60), .D(n59), .Z(n80) );
  AOI22M1P U84 ( .A(transmissionPacket[29]), .B(N103), .C(
        transmissionPacket[28]), .D(N104), .Z(n66) );
  AOI22M1P U85 ( .A(transmissionPacket[27]), .B(N105), .C(
        transmissionPacket[26]), .D(N106), .Z(n65) );
  AOI22M1P U86 ( .A(transmissionPacket[25]), .B(N107), .C(
        transmissionPacket[24]), .D(N108), .Z(n64) );
  AOI22M1P U87 ( .A(transmissionPacket[23]), .B(N109), .C(
        transmissionPacket[22]), .D(N110), .Z(n63) );
  ND4M1P U88 ( .A(n66), .B(n65), .C(n64), .D(n63), .Z(n79) );
  AOI22M1P U89 ( .A(transmissionPacket[20]), .B(N112), .C(
        transmissionPacket[21]), .D(N111), .Z(n70) );
  AOI22M1P U90 ( .A(transmissionPacket[19]), .B(N113), .C(
        transmissionPacket[18]), .D(N114), .Z(n69) );
  AOI22M1P U91 ( .A(transmissionPacket[17]), .B(N115), .C(
        transmissionPacket[16]), .D(N116), .Z(n68) );
  AOI22M1P U92 ( .A(transmissionPacket[15]), .B(N117), .C(
        transmissionPacket[14]), .D(N118), .Z(n67) );
  AND4M1P U93 ( .A(n70), .B(n69), .C(n68), .D(n67), .Z(n77) );
  AOI22M1P U94 ( .A(transmissionPacket[13]), .B(N119), .C(
        transmissionPacket[12]), .D(N120), .Z(n76) );
  AOI22M1P U95 ( .A(transmissionPacket[11]), .B(N121), .C(
        transmissionPacket[10]), .D(N122), .Z(n75) );
  AOI22M1P U96 ( .A(transmissionPacket[9]), .B(N123), .C(transmissionPacket[8]), .D(N124), .Z(n72) );
  AOI22M1P U97 ( .A(transmissionPacket[4]), .B(N128), .C(transmissionPacket[6]), .D(N126), .Z(n71) );
  ND2M1P U98 ( .A(n72), .B(n71), .Z(n73) );
  AOI21M1P U99 ( .A(N125), .B(transmissionPacket[7]), .C(n73), .Z(n74) );
  ND4M1P U100 ( .A(n77), .B(n76), .C(n75), .D(n74), .Z(n78) );
  NR3M1P U101 ( .A(n80), .B(n79), .C(n78), .Z(n83) );
  N1M1P U102 ( .A(n155), .Z(n138) );
  N1M1P U103 ( .A(bitCount[1]), .Z(n128) );
  N1M1P U104 ( .A(bitCount[4]), .Z(n117) );
  ND4DNM1P U105 ( .D(bitCount[3]), .A(n128), .B(n124), .C(n117), .Z(n85) );
  OAI21M1P U106 ( .A(bitCount[0]), .B(n85), .C(bitCount[5]), .Z(n81) );
  AO21CNM1P U107 ( .A(n138), .B(n81), .C(n163), .Z(n82) );
  OAI211M1P U108 ( .A(n83), .B(n131), .C(n153), .D(n82), .Z(N146) );
  N1M1P U109 ( .A(Tx_Ready), .Z(n135) );
  AO21M1P U110 ( .A(n161), .B(n157), .C(n159), .Z(n84) );
  ND3M1P U111 ( .A(Rx_Ready), .B(n135), .C(n84), .Z(n145) );
  N1M1P U112 ( .A(bitCount[5]), .Z(n116) );
  N1M1P U113 ( .A(bitCount[0]), .Z(n130) );
  OR3M1P U114 ( .A(n85), .B(n116), .C(n130), .Z(n86) );
  AOI21M1P U115 ( .A(n135), .B(n86), .C(TxData_Valid), .Z(n143) );
  N1M1P U116 ( .A(transmissionPacket[0]), .Z(n115) );
  AOI22CDNM1P U117 ( .A(TxData[30]), .B(TxData[31]), .C(TxData[31]), .D(
        TxData[30]), .Z(n106) );
  AOI22CDNM1P U118 ( .A(TxData[24]), .B(TxData[25]), .C(TxData[25]), .D(
        TxData[24]), .Z(n90) );
  AOI22CDNM1P U119 ( .A(TxData[26]), .B(TxData[27]), .C(TxData[27]), .D(
        TxData[26]), .Z(n89) );
  N1M1P U120 ( .A(TxData[28]), .Z(n87) );
  AOI22CDNM1P U121 ( .A(TxData[29]), .B(n87), .C(n87), .D(TxData[29]), .Z(n88)
         );
  EN3M1P U122 ( .A(n90), .B(n89), .C(n88), .Z(n105) );
  AOI22CDNM1P U123 ( .A(TxData[6]), .B(TxData[7]), .C(TxData[7]), .D(TxData[6]), .Z(n103) );
  AOI22CDNM1P U124 ( .A(TxData[0]), .B(TxData[1]), .C(TxData[1]), .D(TxData[0]), .Z(n95) );
  AOI22CDNM1P U125 ( .A(TxData[2]), .B(TxData[3]), .C(TxData[3]), .D(TxData[2]), .Z(n94) );
  N1M1P U126 ( .A(TxData[4]), .Z(n91) );
  AOI22CDNM1P U127 ( .A(TxData[5]), .B(n91), .C(n91), .D(TxData[5]), .Z(n92)
         );
  EN3M1P U128 ( .A(n95), .B(n94), .C(n92), .Z(n102) );
  AOI22CDNM1P U129 ( .A(TxData[15]), .B(TxData[16]), .C(TxData[16]), .D(
        TxData[15]), .Z(n99) );
  AOI22CDNM1P U130 ( .A(TxData[17]), .B(TxData[18]), .C(TxData[18]), .D(
        TxData[17]), .Z(n98) );
  N1M1P U131 ( .A(TxData[19]), .Z(n96) );
  AOI22CDNM1P U132 ( .A(TxData[23]), .B(n96), .C(n96), .D(TxData[23]), .Z(n97)
         );
  EN3M1P U133 ( .A(n99), .B(n98), .C(n97), .Z(n100) );
  EN3M1P U134 ( .A(TxData[22]), .B(TxData[14]), .C(n100), .Z(n101) );
  EN3M1P U135 ( .A(n103), .B(n102), .C(n101), .Z(n104) );
  EN3M1P U136 ( .A(n106), .B(n105), .C(n104), .Z(n113) );
  AOI22CDNM1P U137 ( .A(TxData[12]), .B(TxData[13]), .C(TxData[13]), .D(
        TxData[12]), .Z(n109) );
  AOI22CDNM1P U138 ( .A(TxData[8]), .B(TxData[9]), .C(TxData[9]), .D(TxData[8]), .Z(n108) );
  AOI22CDNM1P U139 ( .A(TxData[10]), .B(TxData[11]), .C(TxData[11]), .D(
        TxData[10]), .Z(n107) );
  EN3M1P U140 ( .A(n109), .B(n108), .C(n107), .Z(n110) );
  EN3M1P U141 ( .A(TxData[20]), .B(TxData[21]), .C(n110), .Z(n112) );
  ND2M1P U142 ( .A(n113), .B(n112), .Z(n111) );
  OAI211M1P U143 ( .A(n113), .B(n112), .C(n111), .D(n152), .Z(n114) );
  OAI21M1P U144 ( .A(n152), .B(n115), .C(n114), .Z(n144) );
  NR2M1P U145 ( .A(bitCount[3]), .B(n131), .Z(n121) );
  NR3M1P U146 ( .A(n130), .B(n128), .C(n124), .Z(n120) );
  OAI21M1P U147 ( .A(n120), .B(n131), .C(n153), .Z(n122) );
  NR2M1P U148 ( .A(n121), .B(n122), .Z(n119) );
  ND3M1P U149 ( .A(bitCount[3]), .B(n133), .C(n120), .Z(n118) );
  OAI22M1P U150 ( .A(n119), .B(n116), .C(n117), .D(n118), .Z(n146) );
  AOI22M1P U151 ( .A(bitCount[4]), .B(n119), .C(n118), .D(n117), .Z(n147) );
  AOI22M1P U152 ( .A(bitCount[3]), .B(n122), .C(n121), .D(n120), .Z(n123) );
  N1M1P U153 ( .A(n123), .Z(n148) );
  N1M1P U154 ( .A(n153), .Z(n139) );
  AOI21M1P U155 ( .A(n130), .B(n133), .C(n139), .Z(n129) );
  OA21M1P U156 ( .A(n131), .B(bitCount[1]), .C(n129), .Z(n126) );
  ND3M1P U157 ( .A(bitCount[0]), .B(bitCount[1]), .C(n133), .Z(n125) );
  AOI22M1P U158 ( .A(bitCount[2]), .B(n126), .C(n125), .D(n124), .Z(n149) );
  ND2M1P U159 ( .A(n133), .B(n128), .Z(n127) );
  OAI22M1P U160 ( .A(n129), .B(n128), .C(n130), .D(n127), .Z(n150) );
  AOI22M1P U161 ( .A(bitCount[0]), .B(n153), .C(n131), .D(n130), .Z(n151) );
  N1M1P U162 ( .A(n166), .Z(n141) );
  ND2M1P U163 ( .A(n142), .B(n141), .Z(n154) );
  NR2M1P U164 ( .A(n139), .B(n163), .Z(n132) );
  AOI211M1P U165 ( .A(n138), .B(n139), .C(n133), .D(n132), .Z(n156) );
  NR2M1P U166 ( .A(n161), .B(n145), .Z(n137) );
  N1M1P U167 ( .A(n157), .Z(n134) );
  OR3M1P U168 ( .A(n157), .B(n161), .C(n145), .Z(n136) );
  OAI211M1P U169 ( .A(n137), .B(n134), .C(n135), .D(n136), .Z(n158) );
  AO21CNM1P U170 ( .A(n159), .B(n136), .C(n135), .Z(n160) );
  AO211M1P U171 ( .A(n161), .B(n145), .C(Tx_Ready), .D(n137), .Z(n162) );
  ND3M1P U172 ( .A(n163), .B(n139), .C(n138), .Z(n140) );
endmodule


module tx_2 ( Clk_s, Rst_n, TxData_Valid, TxData, Error_Ack, Rx_Ready, 
        Rx_Error, Tx_Ready, Tx_Error, S_Data );
  input [31:0] TxData;
  input Clk_s, Rst_n, TxData_Valid, Error_Ack, Rx_Ready, Rx_Error;
  output Tx_Ready, Tx_Error, S_Data;
  wire   N100, N101, N102, N103, N104, N105, N106, N107, N108, N109, N110,
         N111, N112, N113, N114, N115, N116, N117, N118, N119, N120, N121,
         N122, N123, N124, N125, N126, N127, N128, N129, N130, N131, N132,
         N146, n17, n18, n19, n20, n21, n22, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167;
  wire   [32:0] transmissionPacket;
  wire   [5:0] bitCount;

  FD4QM1P zeroPatternDetected_reg ( .D(n154), .CP(Clk_s), .SD(Rst_n), .Q(n153)
         );
  FD4QM1P DataTxInProg_reg ( .D(n156), .CP(Clk_s), .SD(Rst_n), .Q(n155) );
  FD4QM1P Tx_Ready_reg ( .D(n143), .CP(Clk_s), .SD(Rst_n), .Q(Tx_Ready) );
  FD2LQM1P \transmissionPacket_reg[1]  ( .D(TxData[0]), .LD(n58), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[1]) );
  FD2LQM1P \transmissionPacket_reg[2]  ( .D(TxData[1]), .LD(n58), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[2]) );
  FD2LQM1P \transmissionPacket_reg[3]  ( .D(TxData[2]), .LD(n58), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[3]) );
  FD2LQM1P \transmissionPacket_reg[4]  ( .D(TxData[3]), .LD(n58), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[4]) );
  FD2LQM1P \transmissionPacket_reg[5]  ( .D(TxData[4]), .LD(n58), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[5]) );
  FD2LQM1P \transmissionPacket_reg[6]  ( .D(TxData[5]), .LD(n58), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[6]) );
  FD2LQM1P \transmissionPacket_reg[7]  ( .D(TxData[6]), .LD(n58), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[7]) );
  FD2LQM1P \transmissionPacket_reg[8]  ( .D(TxData[7]), .LD(n58), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[8]) );
  FD2LQM1P \transmissionPacket_reg[9]  ( .D(TxData[8]), .LD(n58), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[9]) );
  FD2LQM1P \transmissionPacket_reg[10]  ( .D(TxData[9]), .LD(n58), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[10]) );
  FD2LQM1P \transmissionPacket_reg[11]  ( .D(TxData[10]), .LD(n58), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[11]) );
  FD2LQM1P \transmissionPacket_reg[12]  ( .D(TxData[11]), .LD(n58), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[12]) );
  FD2LQM1P \transmissionPacket_reg[13]  ( .D(TxData[12]), .LD(n58), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[13]) );
  FD2LQM1P \transmissionPacket_reg[14]  ( .D(TxData[13]), .LD(n58), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[14]) );
  FD2LQM1P \transmissionPacket_reg[15]  ( .D(TxData[14]), .LD(n58), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[15]) );
  FD2LQM1P \transmissionPacket_reg[16]  ( .D(TxData[15]), .LD(n58), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[16]) );
  FD2LQM1P \transmissionPacket_reg[17]  ( .D(TxData[16]), .LD(n58), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[17]) );
  FD2LQM1P \transmissionPacket_reg[18]  ( .D(TxData[17]), .LD(n58), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[18]) );
  FD2LQM1P \transmissionPacket_reg[19]  ( .D(TxData[18]), .LD(n58), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[19]) );
  FD2LQM1P \transmissionPacket_reg[20]  ( .D(TxData[19]), .LD(n58), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[20]) );
  FD2LQM1P \transmissionPacket_reg[21]  ( .D(TxData[20]), .LD(n58), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[21]) );
  FD2LQM1P \transmissionPacket_reg[22]  ( .D(TxData[21]), .LD(n58), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[22]) );
  FD2LQM1P \transmissionPacket_reg[23]  ( .D(TxData[22]), .LD(n152), .CP(Clk_s), .CD(Rst_n), .Q(transmissionPacket[23]) );
  FD2LQM1P \transmissionPacket_reg[24]  ( .D(TxData[23]), .LD(n152), .CP(Clk_s), .CD(Rst_n), .Q(transmissionPacket[24]) );
  FD2LQM1P \transmissionPacket_reg[25]  ( .D(TxData[24]), .LD(n152), .CP(Clk_s), .CD(Rst_n), .Q(transmissionPacket[25]) );
  FD2LQM1P \transmissionPacket_reg[26]  ( .D(TxData[25]), .LD(n152), .CP(Clk_s), .CD(Rst_n), .Q(transmissionPacket[26]) );
  FD2LQM1P \transmissionPacket_reg[27]  ( .D(TxData[26]), .LD(n152), .CP(Clk_s), .CD(Rst_n), .Q(transmissionPacket[27]) );
  FD2LQM1P \transmissionPacket_reg[28]  ( .D(TxData[27]), .LD(n152), .CP(Clk_s), .CD(Rst_n), .Q(transmissionPacket[28]) );
  FD2LQM1P \transmissionPacket_reg[29]  ( .D(TxData[28]), .LD(n152), .CP(Clk_s), .CD(Rst_n), .Q(transmissionPacket[29]) );
  FD2LQM1P \transmissionPacket_reg[30]  ( .D(TxData[29]), .LD(n152), .CP(Clk_s), .CD(Rst_n), .Q(transmissionPacket[30]) );
  FD2LQM1P \transmissionPacket_reg[31]  ( .D(TxData[30]), .LD(n152), .CP(Clk_s), .CD(Rst_n), .Q(transmissionPacket[31]) );
  FD2LQM1P \transmissionPacket_reg[32]  ( .D(TxData[31]), .LD(n58), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[32]) );
  FD4QM1P \startSequenceCount_reg[1]  ( .D(n158), .CP(Clk_s), .SD(Rst_n), .Q(
        n157) );
  FD4QM1P \startSequenceCount_reg[2]  ( .D(n160), .CP(Clk_s), .SD(Rst_n), .Q(
        n159) );
  FD4QM1P \startSequenceCount_reg[0]  ( .D(n162), .CP(Clk_s), .SD(Rst_n), .Q(
        n161) );
  FD4QM1P startSequence_reg ( .D(n145), .CP(Clk_s), .SD(Rst_n), .Q(n163) );
  FD4QM1P \zeroCount_reg[0]  ( .D(n165), .CP(Clk_s), .SD(Rst_n), .Q(n164) );
  FD4QM1P \zeroCount_reg[1]  ( .D(n167), .CP(Clk_s), .SD(Rst_n), .Q(n166) );
  FD4QM1P S_Data_reg ( .D(N146), .CP(Clk_s), .SD(Rst_n), .Q(S_Data) );
  FD2QM1P \bitCount_reg[0]  ( .D(n151), .CP(Clk_s), .CD(Rst_n), .Q(bitCount[0]) );
  FD2QM1P \bitCount_reg[3]  ( .D(n148), .CP(Clk_s), .CD(Rst_n), .Q(bitCount[3]) );
  FD2QM1P \bitCount_reg[1]  ( .D(n150), .CP(Clk_s), .CD(Rst_n), .Q(bitCount[1]) );
  FD2QM1P \bitCount_reg[5]  ( .D(n146), .CP(Clk_s), .CD(Rst_n), .Q(bitCount[5]) );
  FD2QM1P \bitCount_reg[4]  ( .D(n147), .CP(Clk_s), .CD(Rst_n), .Q(bitCount[4]) );
  FD2QM1P \bitCount_reg[2]  ( .D(n149), .CP(Clk_s), .CD(Rst_n), .Q(bitCount[2]) );
  FD2QM1P \transmissionPacket_reg[0]  ( .D(n144), .CP(Clk_s), .CD(Rst_n), .Q(
        transmissionPacket[0]) );
  ND2BNM1P U3 ( .B(bitCount[1]), .A(bitCount[0]), .Z(n55) );
  ND2BNM1P U4 ( .B(bitCount[0]), .A(bitCount[1]), .Z(n18) );
  N1M1P U5 ( .A(bitCount[2]), .Z(n124) );
  ND4M1P U6 ( .A(n153), .B(n163), .C(n138), .D(n81), .Z(n131) );
  AND2M1P U7 ( .A(Tx_Ready), .B(TxData_Valid), .Z(n152) );
  AOI22DNM1P U8 ( .A(n166), .B(n142), .D(n140), .C(n141), .Z(n17) );
  OA21M1P U9 ( .A(n166), .B(n20), .C(n17), .Z(n167) );
  N1M1P U10 ( .A(n131), .Z(n133) );
  NR2BNM1P U11 ( .B(bitCount[4]), .A(bitCount[5]), .Z(n46) );
  OR2M1P U12 ( .A(bitCount[0]), .B(bitCount[1]), .Z(n54) );
  BUFM2P U13 ( .A(n152), .Z(n58) );
  ND2BNM1P U14 ( .B(n19), .A(n164), .Z(n20) );
  NR2M1P U15 ( .A(n19), .B(n164), .Z(n142) );
  N1M1P U16 ( .A(bitCount[3]), .Z(n57) );
  ND2M1P U17 ( .A(n48), .B(n46), .Z(n43) );
  OA21M1P U18 ( .A(n164), .B(n140), .C(n20), .Z(n165) );
  NR2M1P U19 ( .A(n18), .B(n52), .Z(N106) );
  NR2M1P U20 ( .A(n18), .B(n47), .Z(N130) );
  NR2M1P U21 ( .A(n50), .B(n18), .Z(N102) );
  NR2M1P U22 ( .A(n18), .B(n45), .Z(N126) );
  NR2M1P U23 ( .A(n18), .B(n44), .Z(N122) );
  NR2M1P U24 ( .A(n18), .B(n43), .Z(N118) );
  NR2M1P U25 ( .A(n18), .B(n42), .Z(N114) );
  NR2M1P U26 ( .A(n56), .B(n18), .Z(N110) );
  ND2M1P U27 ( .A(n41), .B(n40), .Z(n19) );
  AOI22M1P U28 ( .A(transmissionPacket[13]), .B(N119), .C(
        transmissionPacket[12]), .D(N120), .Z(n21) );
  AOI22M1P U29 ( .A(transmissionPacket[22]), .B(N110), .C(
        transmissionPacket[21]), .D(N111), .Z(n22) );
  AOI22M1P U30 ( .A(transmissionPacket[23]), .B(N109), .C(
        transmissionPacket[20]), .D(N112), .Z(n29) );
  AOI22M1P U31 ( .A(transmissionPacket[2]), .B(N130), .C(transmissionPacket[1]), .D(N131), .Z(n30) );
  AOI22M1P U32 ( .A(transmissionPacket[4]), .B(N128), .C(transmissionPacket[6]), .D(N126), .Z(n31) );
  AOI22M1P U33 ( .A(transmissionPacket[5]), .B(N127), .C(transmissionPacket[3]), .D(N129), .Z(n32) );
  AOI22M1P U34 ( .A(transmissionPacket[7]), .B(N125), .C(transmissionPacket[9]), .D(N123), .Z(n33) );
  AOI22M1P U35 ( .A(transmissionPacket[11]), .B(N121), .C(
        transmissionPacket[10]), .D(N122), .Z(n34) );
  ND4M1P U36 ( .A(n69), .B(n68), .C(n67), .D(n21), .Z(n35) );
  ND4M1P U37 ( .A(n65), .B(n64), .C(n29), .D(n22), .Z(n36) );
  ND4M1P U38 ( .A(n30), .B(n60), .C(n59), .D(n66), .Z(n37) );
  ND4M1P U39 ( .A(n34), .B(n33), .C(n32), .D(n31), .Z(n38) );
  ND3M1P U40 ( .A(n138), .B(n153), .C(n163), .Z(n39) );
  NR3M1P U41 ( .A(n37), .B(n36), .C(n35), .Z(n40) );
  AOI211M1P U42 ( .A(N124), .B(transmissionPacket[8]), .C(n39), .D(n38), .Z(
        n41) );
  NR2M1P U43 ( .A(n54), .B(n50), .Z(N100) );
  NR2M1P U44 ( .A(n56), .B(n53), .Z(N111) );
  NR2M1P U45 ( .A(n54), .B(n42), .Z(N112) );
  NR2M1P U46 ( .A(n42), .B(n55), .Z(N113) );
  NR2M1P U47 ( .A(n53), .B(n42), .Z(N115) );
  NR2M1P U48 ( .A(n54), .B(n43), .Z(N116) );
  NR2M1P U49 ( .A(n55), .B(n43), .Z(N117) );
  NR2M1P U50 ( .A(n53), .B(n43), .Z(N119) );
  NR2M1P U51 ( .A(n50), .B(n55), .Z(N101) );
  NR2M1P U52 ( .A(n54), .B(n44), .Z(N120) );
  NR2M1P U53 ( .A(n55), .B(n44), .Z(N121) );
  NR2M1P U54 ( .A(n53), .B(n44), .Z(N123) );
  NR2M1P U55 ( .A(n54), .B(n45), .Z(N124) );
  NR2M1P U56 ( .A(n55), .B(n45), .Z(N125) );
  NR2M1P U57 ( .A(n53), .B(n45), .Z(N127) );
  NR2M1P U58 ( .A(n54), .B(n47), .Z(N128) );
  NR2M1P U59 ( .A(n55), .B(n47), .Z(N129) );
  NR2M1P U60 ( .A(n53), .B(n47), .Z(N131) );
  NR3M1P U61 ( .A(bitCount[4]), .B(n54), .C(n49), .Z(N132) );
  NR2M1P U62 ( .A(n50), .B(n53), .Z(N103) );
  NR2M1P U63 ( .A(n54), .B(n52), .Z(N104) );
  NR2M1P U64 ( .A(n55), .B(n52), .Z(N105) );
  NR2M1P U65 ( .A(n53), .B(n52), .Z(N107) );
  NR2M1P U66 ( .A(n54), .B(n56), .Z(N108) );
  NR2M1P U67 ( .A(n56), .B(n55), .Z(N109) );
  NR2M1P U68 ( .A(bitCount[5]), .B(bitCount[4]), .Z(n51) );
  NR2M1P U69 ( .A(bitCount[2]), .B(bitCount[3]), .Z(n48) );
  ND2M1P U70 ( .A(n51), .B(n48), .Z(n50) );
  ND3M1P U71 ( .A(n51), .B(bitCount[3]), .C(n124), .Z(n56) );
  ND2M1P U72 ( .A(bitCount[1]), .B(bitCount[0]), .Z(n53) );
  ND3M1P U73 ( .A(n51), .B(bitCount[2]), .C(bitCount[3]), .Z(n42) );
  ND3M1P U74 ( .A(bitCount[2]), .B(n46), .C(n57), .Z(n44) );
  ND3M1P U75 ( .A(bitCount[3]), .B(n46), .C(n124), .Z(n45) );
  ND3M1P U76 ( .A(bitCount[2]), .B(bitCount[3]), .C(n46), .Z(n47) );
  ND2M1P U77 ( .A(bitCount[5]), .B(n48), .Z(n49) );
  ND3M1P U78 ( .A(bitCount[2]), .B(n51), .C(n57), .Z(n52) );
  AOI22M1P U79 ( .A(transmissionPacket[5]), .B(N127), .C(transmissionPacket[3]), .D(N129), .Z(n62) );
  AOI22M1P U80 ( .A(transmissionPacket[2]), .B(N130), .C(transmissionPacket[1]), .D(N131), .Z(n61) );
  AOI22M1P U81 ( .A(transmissionPacket[32]), .B(N100), .C(
        transmissionPacket[0]), .D(N132), .Z(n60) );
  AOI22M1P U82 ( .A(transmissionPacket[30]), .B(N102), .C(
        transmissionPacket[31]), .D(N101), .Z(n59) );
  ND4M1P U83 ( .A(n62), .B(n61), .C(n60), .D(n59), .Z(n80) );
  AOI22M1P U84 ( .A(transmissionPacket[29]), .B(N103), .C(
        transmissionPacket[28]), .D(N104), .Z(n66) );
  AOI22M1P U85 ( .A(transmissionPacket[27]), .B(N105), .C(
        transmissionPacket[26]), .D(N106), .Z(n65) );
  AOI22M1P U86 ( .A(transmissionPacket[25]), .B(N107), .C(
        transmissionPacket[24]), .D(N108), .Z(n64) );
  AOI22M1P U87 ( .A(transmissionPacket[23]), .B(N109), .C(
        transmissionPacket[22]), .D(N110), .Z(n63) );
  ND4M1P U88 ( .A(n66), .B(n65), .C(n64), .D(n63), .Z(n79) );
  AOI22M1P U89 ( .A(transmissionPacket[20]), .B(N112), .C(
        transmissionPacket[21]), .D(N111), .Z(n70) );
  AOI22M1P U90 ( .A(transmissionPacket[19]), .B(N113), .C(
        transmissionPacket[18]), .D(N114), .Z(n69) );
  AOI22M1P U91 ( .A(transmissionPacket[17]), .B(N115), .C(
        transmissionPacket[16]), .D(N116), .Z(n68) );
  AOI22M1P U92 ( .A(transmissionPacket[15]), .B(N117), .C(
        transmissionPacket[14]), .D(N118), .Z(n67) );
  AND4M1P U93 ( .A(n70), .B(n69), .C(n68), .D(n67), .Z(n77) );
  AOI22M1P U94 ( .A(transmissionPacket[13]), .B(N119), .C(
        transmissionPacket[12]), .D(N120), .Z(n76) );
  AOI22M1P U95 ( .A(transmissionPacket[11]), .B(N121), .C(
        transmissionPacket[10]), .D(N122), .Z(n75) );
  AOI22M1P U96 ( .A(transmissionPacket[9]), .B(N123), .C(transmissionPacket[8]), .D(N124), .Z(n72) );
  AOI22M1P U97 ( .A(transmissionPacket[4]), .B(N128), .C(transmissionPacket[6]), .D(N126), .Z(n71) );
  ND2M1P U98 ( .A(n72), .B(n71), .Z(n73) );
  AOI21M1P U99 ( .A(N125), .B(transmissionPacket[7]), .C(n73), .Z(n74) );
  ND4M1P U100 ( .A(n77), .B(n76), .C(n75), .D(n74), .Z(n78) );
  NR3M1P U101 ( .A(n80), .B(n79), .C(n78), .Z(n83) );
  N1M1P U102 ( .A(n155), .Z(n138) );
  N1M1P U103 ( .A(bitCount[1]), .Z(n128) );
  N1M1P U104 ( .A(bitCount[4]), .Z(n117) );
  ND4DNM1P U105 ( .D(bitCount[3]), .A(n128), .B(n124), .C(n117), .Z(n85) );
  OAI21M1P U106 ( .A(bitCount[0]), .B(n85), .C(bitCount[5]), .Z(n81) );
  AO21CNM1P U107 ( .A(n138), .B(n81), .C(n163), .Z(n82) );
  OAI211M1P U108 ( .A(n83), .B(n131), .C(n153), .D(n82), .Z(N146) );
  N1M1P U109 ( .A(Tx_Ready), .Z(n135) );
  AO21M1P U110 ( .A(n161), .B(n157), .C(n159), .Z(n84) );
  ND3M1P U111 ( .A(Rx_Ready), .B(n135), .C(n84), .Z(n145) );
  N1M1P U112 ( .A(bitCount[5]), .Z(n116) );
  N1M1P U113 ( .A(bitCount[0]), .Z(n130) );
  OR3M1P U114 ( .A(n85), .B(n116), .C(n130), .Z(n86) );
  AOI21M1P U115 ( .A(n135), .B(n86), .C(TxData_Valid), .Z(n143) );
  N1M1P U116 ( .A(transmissionPacket[0]), .Z(n115) );
  AOI22CDNM1P U117 ( .A(TxData[30]), .B(TxData[31]), .C(TxData[31]), .D(
        TxData[30]), .Z(n106) );
  AOI22CDNM1P U118 ( .A(TxData[24]), .B(TxData[25]), .C(TxData[25]), .D(
        TxData[24]), .Z(n90) );
  AOI22CDNM1P U119 ( .A(TxData[26]), .B(TxData[27]), .C(TxData[27]), .D(
        TxData[26]), .Z(n89) );
  N1M1P U120 ( .A(TxData[28]), .Z(n87) );
  AOI22CDNM1P U121 ( .A(TxData[29]), .B(n87), .C(n87), .D(TxData[29]), .Z(n88)
         );
  EN3M1P U122 ( .A(n90), .B(n89), .C(n88), .Z(n105) );
  AOI22CDNM1P U123 ( .A(TxData[6]), .B(TxData[7]), .C(TxData[7]), .D(TxData[6]), .Z(n103) );
  AOI22CDNM1P U124 ( .A(TxData[0]), .B(TxData[1]), .C(TxData[1]), .D(TxData[0]), .Z(n95) );
  AOI22CDNM1P U125 ( .A(TxData[2]), .B(TxData[3]), .C(TxData[3]), .D(TxData[2]), .Z(n94) );
  N1M1P U126 ( .A(TxData[4]), .Z(n91) );
  AOI22CDNM1P U127 ( .A(TxData[5]), .B(n91), .C(n91), .D(TxData[5]), .Z(n92)
         );
  EN3M1P U128 ( .A(n95), .B(n94), .C(n92), .Z(n102) );
  AOI22CDNM1P U129 ( .A(TxData[15]), .B(TxData[16]), .C(TxData[16]), .D(
        TxData[15]), .Z(n99) );
  AOI22CDNM1P U130 ( .A(TxData[17]), .B(TxData[18]), .C(TxData[18]), .D(
        TxData[17]), .Z(n98) );
  N1M1P U131 ( .A(TxData[19]), .Z(n96) );
  AOI22CDNM1P U132 ( .A(TxData[23]), .B(n96), .C(n96), .D(TxData[23]), .Z(n97)
         );
  EN3M1P U133 ( .A(n99), .B(n98), .C(n97), .Z(n100) );
  EN3M1P U134 ( .A(TxData[22]), .B(TxData[14]), .C(n100), .Z(n101) );
  EN3M1P U135 ( .A(n103), .B(n102), .C(n101), .Z(n104) );
  EN3M1P U136 ( .A(n106), .B(n105), .C(n104), .Z(n113) );
  AOI22CDNM1P U137 ( .A(TxData[12]), .B(TxData[13]), .C(TxData[13]), .D(
        TxData[12]), .Z(n109) );
  AOI22CDNM1P U138 ( .A(TxData[8]), .B(TxData[9]), .C(TxData[9]), .D(TxData[8]), .Z(n108) );
  AOI22CDNM1P U139 ( .A(TxData[10]), .B(TxData[11]), .C(TxData[11]), .D(
        TxData[10]), .Z(n107) );
  EN3M1P U140 ( .A(n109), .B(n108), .C(n107), .Z(n110) );
  EN3M1P U141 ( .A(TxData[20]), .B(TxData[21]), .C(n110), .Z(n112) );
  ND2M1P U142 ( .A(n113), .B(n112), .Z(n111) );
  OAI211M1P U143 ( .A(n113), .B(n112), .C(n111), .D(n152), .Z(n114) );
  OAI21M1P U144 ( .A(n152), .B(n115), .C(n114), .Z(n144) );
  NR2M1P U145 ( .A(bitCount[3]), .B(n131), .Z(n121) );
  NR3M1P U146 ( .A(n130), .B(n128), .C(n124), .Z(n120) );
  OAI21M1P U147 ( .A(n120), .B(n131), .C(n153), .Z(n122) );
  NR2M1P U148 ( .A(n121), .B(n122), .Z(n119) );
  ND3M1P U149 ( .A(bitCount[3]), .B(n133), .C(n120), .Z(n118) );
  OAI22M1P U150 ( .A(n119), .B(n116), .C(n117), .D(n118), .Z(n146) );
  AOI22M1P U151 ( .A(bitCount[4]), .B(n119), .C(n118), .D(n117), .Z(n147) );
  AOI22M1P U152 ( .A(bitCount[3]), .B(n122), .C(n121), .D(n120), .Z(n123) );
  N1M1P U153 ( .A(n123), .Z(n148) );
  N1M1P U154 ( .A(n153), .Z(n139) );
  AOI21M1P U155 ( .A(n130), .B(n133), .C(n139), .Z(n129) );
  OA21M1P U156 ( .A(n131), .B(bitCount[1]), .C(n129), .Z(n126) );
  ND3M1P U157 ( .A(bitCount[0]), .B(bitCount[1]), .C(n133), .Z(n125) );
  AOI22M1P U158 ( .A(bitCount[2]), .B(n126), .C(n125), .D(n124), .Z(n149) );
  ND2M1P U159 ( .A(n133), .B(n128), .Z(n127) );
  OAI22M1P U160 ( .A(n129), .B(n128), .C(n130), .D(n127), .Z(n150) );
  AOI22M1P U161 ( .A(bitCount[0]), .B(n153), .C(n131), .D(n130), .Z(n151) );
  N1M1P U162 ( .A(n166), .Z(n141) );
  ND2M1P U163 ( .A(n142), .B(n141), .Z(n154) );
  NR2M1P U164 ( .A(n139), .B(n163), .Z(n132) );
  AOI211M1P U165 ( .A(n138), .B(n139), .C(n133), .D(n132), .Z(n156) );
  NR2M1P U166 ( .A(n161), .B(n145), .Z(n137) );
  N1M1P U167 ( .A(n157), .Z(n134) );
  OR3M1P U168 ( .A(n157), .B(n161), .C(n145), .Z(n136) );
  OAI211M1P U169 ( .A(n137), .B(n134), .C(n135), .D(n136), .Z(n158) );
  AO21CNM1P U170 ( .A(n159), .B(n136), .C(n135), .Z(n160) );
  AO211M1P U171 ( .A(n161), .B(n145), .C(Tx_Ready), .D(n137), .Z(n162) );
  ND3M1P U172 ( .A(n163), .B(n139), .C(n138), .Z(n140) );
endmodule


module tx_3 ( Clk_s, Rst_n, TxData_Valid, TxData, Error_Ack, Rx_Ready, 
        Rx_Error, Tx_Ready, Tx_Error, S_Data );
  input [31:0] TxData;
  input Clk_s, Rst_n, TxData_Valid, Error_Ack, Rx_Ready, Rx_Error;
  output Tx_Ready, Tx_Error, S_Data;
  wire   N100, N101, N102, N103, N104, N105, N106, N107, N108, N109, N110,
         N111, N112, N113, N114, N115, N116, N117, N118, N119, N120, N121,
         N122, N123, N124, N125, N126, N127, N128, N129, N130, N131, N132,
         N146, n17, n18, n19, n20, n21, n22, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167;
  wire   [32:0] transmissionPacket;
  wire   [5:0] bitCount;

  FD4QM1P zeroPatternDetected_reg ( .D(n154), .CP(Clk_s), .SD(Rst_n), .Q(n153)
         );
  FD4QM1P DataTxInProg_reg ( .D(n156), .CP(Clk_s), .SD(Rst_n), .Q(n155) );
  FD4QM1P Tx_Ready_reg ( .D(n143), .CP(Clk_s), .SD(Rst_n), .Q(Tx_Ready) );
  FD2LQM1P \transmissionPacket_reg[1]  ( .D(TxData[0]), .LD(n58), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[1]) );
  FD2LQM1P \transmissionPacket_reg[2]  ( .D(TxData[1]), .LD(n58), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[2]) );
  FD2LQM1P \transmissionPacket_reg[3]  ( .D(TxData[2]), .LD(n58), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[3]) );
  FD2LQM1P \transmissionPacket_reg[4]  ( .D(TxData[3]), .LD(n58), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[4]) );
  FD2LQM1P \transmissionPacket_reg[5]  ( .D(TxData[4]), .LD(n58), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[5]) );
  FD2LQM1P \transmissionPacket_reg[6]  ( .D(TxData[5]), .LD(n58), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[6]) );
  FD2LQM1P \transmissionPacket_reg[7]  ( .D(TxData[6]), .LD(n58), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[7]) );
  FD2LQM1P \transmissionPacket_reg[8]  ( .D(TxData[7]), .LD(n58), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[8]) );
  FD2LQM1P \transmissionPacket_reg[9]  ( .D(TxData[8]), .LD(n58), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[9]) );
  FD2LQM1P \transmissionPacket_reg[10]  ( .D(TxData[9]), .LD(n58), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[10]) );
  FD2LQM1P \transmissionPacket_reg[11]  ( .D(TxData[10]), .LD(n58), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[11]) );
  FD2LQM1P \transmissionPacket_reg[12]  ( .D(TxData[11]), .LD(n58), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[12]) );
  FD2LQM1P \transmissionPacket_reg[13]  ( .D(TxData[12]), .LD(n58), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[13]) );
  FD2LQM1P \transmissionPacket_reg[14]  ( .D(TxData[13]), .LD(n58), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[14]) );
  FD2LQM1P \transmissionPacket_reg[15]  ( .D(TxData[14]), .LD(n58), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[15]) );
  FD2LQM1P \transmissionPacket_reg[16]  ( .D(TxData[15]), .LD(n58), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[16]) );
  FD2LQM1P \transmissionPacket_reg[17]  ( .D(TxData[16]), .LD(n58), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[17]) );
  FD2LQM1P \transmissionPacket_reg[18]  ( .D(TxData[17]), .LD(n58), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[18]) );
  FD2LQM1P \transmissionPacket_reg[19]  ( .D(TxData[18]), .LD(n58), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[19]) );
  FD2LQM1P \transmissionPacket_reg[20]  ( .D(TxData[19]), .LD(n58), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[20]) );
  FD2LQM1P \transmissionPacket_reg[21]  ( .D(TxData[20]), .LD(n58), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[21]) );
  FD2LQM1P \transmissionPacket_reg[22]  ( .D(TxData[21]), .LD(n58), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[22]) );
  FD2LQM1P \transmissionPacket_reg[23]  ( .D(TxData[22]), .LD(n152), .CP(Clk_s), .CD(Rst_n), .Q(transmissionPacket[23]) );
  FD2LQM1P \transmissionPacket_reg[24]  ( .D(TxData[23]), .LD(n152), .CP(Clk_s), .CD(Rst_n), .Q(transmissionPacket[24]) );
  FD2LQM1P \transmissionPacket_reg[25]  ( .D(TxData[24]), .LD(n152), .CP(Clk_s), .CD(Rst_n), .Q(transmissionPacket[25]) );
  FD2LQM1P \transmissionPacket_reg[26]  ( .D(TxData[25]), .LD(n152), .CP(Clk_s), .CD(Rst_n), .Q(transmissionPacket[26]) );
  FD2LQM1P \transmissionPacket_reg[27]  ( .D(TxData[26]), .LD(n152), .CP(Clk_s), .CD(Rst_n), .Q(transmissionPacket[27]) );
  FD2LQM1P \transmissionPacket_reg[28]  ( .D(TxData[27]), .LD(n152), .CP(Clk_s), .CD(Rst_n), .Q(transmissionPacket[28]) );
  FD2LQM1P \transmissionPacket_reg[29]  ( .D(TxData[28]), .LD(n152), .CP(Clk_s), .CD(Rst_n), .Q(transmissionPacket[29]) );
  FD2LQM1P \transmissionPacket_reg[30]  ( .D(TxData[29]), .LD(n152), .CP(Clk_s), .CD(Rst_n), .Q(transmissionPacket[30]) );
  FD2LQM1P \transmissionPacket_reg[31]  ( .D(TxData[30]), .LD(n152), .CP(Clk_s), .CD(Rst_n), .Q(transmissionPacket[31]) );
  FD2LQM1P \transmissionPacket_reg[32]  ( .D(TxData[31]), .LD(n58), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[32]) );
  FD4QM1P \startSequenceCount_reg[1]  ( .D(n158), .CP(Clk_s), .SD(Rst_n), .Q(
        n157) );
  FD4QM1P \startSequenceCount_reg[2]  ( .D(n160), .CP(Clk_s), .SD(Rst_n), .Q(
        n159) );
  FD4QM1P \startSequenceCount_reg[0]  ( .D(n162), .CP(Clk_s), .SD(Rst_n), .Q(
        n161) );
  FD4QM1P startSequence_reg ( .D(n145), .CP(Clk_s), .SD(Rst_n), .Q(n163) );
  FD4QM1P \zeroCount_reg[0]  ( .D(n165), .CP(Clk_s), .SD(Rst_n), .Q(n164) );
  FD4QM1P \zeroCount_reg[1]  ( .D(n167), .CP(Clk_s), .SD(Rst_n), .Q(n166) );
  FD4QM1P S_Data_reg ( .D(N146), .CP(Clk_s), .SD(Rst_n), .Q(S_Data) );
  FD2QM1P \bitCount_reg[0]  ( .D(n151), .CP(Clk_s), .CD(Rst_n), .Q(bitCount[0]) );
  FD2QM1P \bitCount_reg[3]  ( .D(n148), .CP(Clk_s), .CD(Rst_n), .Q(bitCount[3]) );
  FD2QM1P \bitCount_reg[1]  ( .D(n150), .CP(Clk_s), .CD(Rst_n), .Q(bitCount[1]) );
  FD2QM1P \bitCount_reg[5]  ( .D(n146), .CP(Clk_s), .CD(Rst_n), .Q(bitCount[5]) );
  FD2QM1P \bitCount_reg[4]  ( .D(n147), .CP(Clk_s), .CD(Rst_n), .Q(bitCount[4]) );
  FD2QM1P \bitCount_reg[2]  ( .D(n149), .CP(Clk_s), .CD(Rst_n), .Q(bitCount[2]) );
  FD2QM1P \transmissionPacket_reg[0]  ( .D(n144), .CP(Clk_s), .CD(Rst_n), .Q(
        transmissionPacket[0]) );
  ND2BNM1P U3 ( .B(bitCount[0]), .A(bitCount[1]), .Z(n18) );
  ND2BNM1P U4 ( .B(bitCount[1]), .A(bitCount[0]), .Z(n55) );
  OR2M1P U5 ( .A(bitCount[0]), .B(bitCount[1]), .Z(n54) );
  ND2M1P U6 ( .A(bitCount[1]), .B(bitCount[0]), .Z(n53) );
  N1M1P U7 ( .A(bitCount[2]), .Z(n124) );
  ND4M1P U8 ( .A(n153), .B(n163), .C(n138), .D(n81), .Z(n131) );
  AND2M1P U9 ( .A(Tx_Ready), .B(TxData_Valid), .Z(n152) );
  AOI22DNM1P U10 ( .A(n166), .B(n142), .D(n140), .C(n141), .Z(n17) );
  OA21M1P U11 ( .A(n166), .B(n20), .C(n17), .Z(n167) );
  N1M1P U12 ( .A(n131), .Z(n133) );
  NR2BNM1P U13 ( .B(bitCount[4]), .A(bitCount[5]), .Z(n46) );
  BUFM2P U14 ( .A(n152), .Z(n58) );
  ND2BNM1P U15 ( .B(n19), .A(n164), .Z(n20) );
  NR2M1P U16 ( .A(n19), .B(n164), .Z(n142) );
  N1M1P U17 ( .A(bitCount[3]), .Z(n57) );
  ND2M1P U18 ( .A(n48), .B(n46), .Z(n43) );
  OA21M1P U19 ( .A(n164), .B(n140), .C(n20), .Z(n165) );
  NR2M1P U20 ( .A(n18), .B(n52), .Z(N106) );
  NR2M1P U21 ( .A(n18), .B(n47), .Z(N130) );
  NR2M1P U22 ( .A(n50), .B(n18), .Z(N102) );
  NR2M1P U23 ( .A(n18), .B(n45), .Z(N126) );
  NR2M1P U24 ( .A(n18), .B(n44), .Z(N122) );
  NR2M1P U25 ( .A(n18), .B(n43), .Z(N118) );
  NR2M1P U26 ( .A(n18), .B(n42), .Z(N114) );
  NR2M1P U27 ( .A(n56), .B(n18), .Z(N110) );
  ND2M1P U28 ( .A(n41), .B(n40), .Z(n19) );
  AOI22M1P U29 ( .A(transmissionPacket[13]), .B(N119), .C(
        transmissionPacket[12]), .D(N120), .Z(n21) );
  AOI22M1P U30 ( .A(transmissionPacket[22]), .B(N110), .C(
        transmissionPacket[21]), .D(N111), .Z(n22) );
  AOI22M1P U31 ( .A(transmissionPacket[23]), .B(N109), .C(
        transmissionPacket[20]), .D(N112), .Z(n29) );
  AOI22M1P U32 ( .A(transmissionPacket[2]), .B(N130), .C(transmissionPacket[1]), .D(N131), .Z(n30) );
  AOI22M1P U33 ( .A(transmissionPacket[4]), .B(N128), .C(transmissionPacket[6]), .D(N126), .Z(n31) );
  AOI22M1P U34 ( .A(transmissionPacket[5]), .B(N127), .C(transmissionPacket[3]), .D(N129), .Z(n32) );
  AOI22M1P U35 ( .A(transmissionPacket[7]), .B(N125), .C(transmissionPacket[9]), .D(N123), .Z(n33) );
  AOI22M1P U36 ( .A(transmissionPacket[11]), .B(N121), .C(
        transmissionPacket[10]), .D(N122), .Z(n34) );
  ND4M1P U37 ( .A(n69), .B(n68), .C(n67), .D(n21), .Z(n35) );
  ND4M1P U38 ( .A(n65), .B(n64), .C(n29), .D(n22), .Z(n36) );
  ND4M1P U39 ( .A(n30), .B(n60), .C(n59), .D(n66), .Z(n37) );
  ND4M1P U40 ( .A(n34), .B(n33), .C(n32), .D(n31), .Z(n38) );
  ND3M1P U41 ( .A(n138), .B(n153), .C(n163), .Z(n39) );
  NR3M1P U42 ( .A(n37), .B(n36), .C(n35), .Z(n40) );
  AOI211M1P U43 ( .A(N124), .B(transmissionPacket[8]), .C(n39), .D(n38), .Z(
        n41) );
  NR2M1P U44 ( .A(n54), .B(n50), .Z(N100) );
  NR2M1P U45 ( .A(n56), .B(n53), .Z(N111) );
  NR2M1P U46 ( .A(n54), .B(n42), .Z(N112) );
  NR2M1P U47 ( .A(n42), .B(n55), .Z(N113) );
  NR2M1P U48 ( .A(n53), .B(n42), .Z(N115) );
  NR2M1P U49 ( .A(n54), .B(n43), .Z(N116) );
  NR2M1P U50 ( .A(n55), .B(n43), .Z(N117) );
  NR2M1P U51 ( .A(n53), .B(n43), .Z(N119) );
  NR2M1P U52 ( .A(n50), .B(n55), .Z(N101) );
  NR2M1P U53 ( .A(n54), .B(n44), .Z(N120) );
  NR2M1P U54 ( .A(n55), .B(n44), .Z(N121) );
  NR2M1P U55 ( .A(n53), .B(n44), .Z(N123) );
  NR2M1P U56 ( .A(n54), .B(n45), .Z(N124) );
  NR2M1P U57 ( .A(n55), .B(n45), .Z(N125) );
  NR2M1P U58 ( .A(n53), .B(n45), .Z(N127) );
  NR2M1P U59 ( .A(n54), .B(n47), .Z(N128) );
  NR2M1P U60 ( .A(n55), .B(n47), .Z(N129) );
  NR2M1P U61 ( .A(n53), .B(n47), .Z(N131) );
  NR3M1P U62 ( .A(bitCount[4]), .B(n54), .C(n49), .Z(N132) );
  NR2M1P U63 ( .A(n50), .B(n53), .Z(N103) );
  NR2M1P U64 ( .A(n54), .B(n52), .Z(N104) );
  NR2M1P U65 ( .A(n55), .B(n52), .Z(N105) );
  NR2M1P U66 ( .A(n53), .B(n52), .Z(N107) );
  NR2M1P U67 ( .A(n54), .B(n56), .Z(N108) );
  NR2M1P U68 ( .A(n56), .B(n55), .Z(N109) );
  NR2M1P U69 ( .A(bitCount[5]), .B(bitCount[4]), .Z(n51) );
  NR2M1P U70 ( .A(bitCount[2]), .B(bitCount[3]), .Z(n48) );
  ND2M1P U71 ( .A(n51), .B(n48), .Z(n50) );
  ND3M1P U72 ( .A(n51), .B(bitCount[3]), .C(n124), .Z(n56) );
  ND3M1P U73 ( .A(n51), .B(bitCount[2]), .C(bitCount[3]), .Z(n42) );
  ND3M1P U74 ( .A(bitCount[2]), .B(n46), .C(n57), .Z(n44) );
  ND3M1P U75 ( .A(bitCount[3]), .B(n46), .C(n124), .Z(n45) );
  ND3M1P U76 ( .A(bitCount[2]), .B(bitCount[3]), .C(n46), .Z(n47) );
  ND2M1P U77 ( .A(bitCount[5]), .B(n48), .Z(n49) );
  ND3M1P U78 ( .A(bitCount[2]), .B(n51), .C(n57), .Z(n52) );
  AOI22M1P U79 ( .A(transmissionPacket[5]), .B(N127), .C(transmissionPacket[3]), .D(N129), .Z(n62) );
  AOI22M1P U80 ( .A(transmissionPacket[2]), .B(N130), .C(transmissionPacket[1]), .D(N131), .Z(n61) );
  AOI22M1P U81 ( .A(transmissionPacket[32]), .B(N100), .C(
        transmissionPacket[0]), .D(N132), .Z(n60) );
  AOI22M1P U82 ( .A(transmissionPacket[30]), .B(N102), .C(
        transmissionPacket[31]), .D(N101), .Z(n59) );
  ND4M1P U83 ( .A(n62), .B(n61), .C(n60), .D(n59), .Z(n80) );
  AOI22M1P U84 ( .A(transmissionPacket[29]), .B(N103), .C(
        transmissionPacket[28]), .D(N104), .Z(n66) );
  AOI22M1P U85 ( .A(transmissionPacket[27]), .B(N105), .C(
        transmissionPacket[26]), .D(N106), .Z(n65) );
  AOI22M1P U86 ( .A(transmissionPacket[25]), .B(N107), .C(
        transmissionPacket[24]), .D(N108), .Z(n64) );
  AOI22M1P U87 ( .A(transmissionPacket[23]), .B(N109), .C(
        transmissionPacket[22]), .D(N110), .Z(n63) );
  ND4M1P U88 ( .A(n66), .B(n65), .C(n64), .D(n63), .Z(n79) );
  AOI22M1P U89 ( .A(transmissionPacket[20]), .B(N112), .C(
        transmissionPacket[21]), .D(N111), .Z(n70) );
  AOI22M1P U90 ( .A(transmissionPacket[19]), .B(N113), .C(
        transmissionPacket[18]), .D(N114), .Z(n69) );
  AOI22M1P U91 ( .A(transmissionPacket[17]), .B(N115), .C(
        transmissionPacket[16]), .D(N116), .Z(n68) );
  AOI22M1P U92 ( .A(transmissionPacket[15]), .B(N117), .C(
        transmissionPacket[14]), .D(N118), .Z(n67) );
  AND4M1P U93 ( .A(n70), .B(n69), .C(n68), .D(n67), .Z(n77) );
  AOI22M1P U94 ( .A(transmissionPacket[13]), .B(N119), .C(
        transmissionPacket[12]), .D(N120), .Z(n76) );
  AOI22M1P U95 ( .A(transmissionPacket[11]), .B(N121), .C(
        transmissionPacket[10]), .D(N122), .Z(n75) );
  AOI22M1P U96 ( .A(transmissionPacket[9]), .B(N123), .C(transmissionPacket[8]), .D(N124), .Z(n72) );
  AOI22M1P U97 ( .A(transmissionPacket[4]), .B(N128), .C(transmissionPacket[6]), .D(N126), .Z(n71) );
  ND2M1P U98 ( .A(n72), .B(n71), .Z(n73) );
  AOI21M1P U99 ( .A(N125), .B(transmissionPacket[7]), .C(n73), .Z(n74) );
  ND4M1P U100 ( .A(n77), .B(n76), .C(n75), .D(n74), .Z(n78) );
  NR3M1P U101 ( .A(n80), .B(n79), .C(n78), .Z(n83) );
  N1M1P U102 ( .A(n155), .Z(n138) );
  N1M1P U103 ( .A(bitCount[1]), .Z(n128) );
  N1M1P U104 ( .A(bitCount[4]), .Z(n117) );
  ND4DNM1P U105 ( .D(bitCount[3]), .A(n128), .B(n124), .C(n117), .Z(n85) );
  OAI21M1P U106 ( .A(bitCount[0]), .B(n85), .C(bitCount[5]), .Z(n81) );
  AO21CNM1P U107 ( .A(n138), .B(n81), .C(n163), .Z(n82) );
  OAI211M1P U108 ( .A(n83), .B(n131), .C(n153), .D(n82), .Z(N146) );
  N1M1P U109 ( .A(Tx_Ready), .Z(n135) );
  AO21M1P U110 ( .A(n161), .B(n157), .C(n159), .Z(n84) );
  ND3M1P U111 ( .A(Rx_Ready), .B(n135), .C(n84), .Z(n145) );
  N1M1P U112 ( .A(bitCount[5]), .Z(n116) );
  N1M1P U113 ( .A(bitCount[0]), .Z(n130) );
  OR3M1P U114 ( .A(n85), .B(n116), .C(n130), .Z(n86) );
  AOI21M1P U115 ( .A(n135), .B(n86), .C(TxData_Valid), .Z(n143) );
  N1M1P U116 ( .A(transmissionPacket[0]), .Z(n115) );
  AOI22CDNM1P U117 ( .A(TxData[30]), .B(TxData[31]), .C(TxData[31]), .D(
        TxData[30]), .Z(n106) );
  AOI22CDNM1P U118 ( .A(TxData[24]), .B(TxData[25]), .C(TxData[25]), .D(
        TxData[24]), .Z(n90) );
  AOI22CDNM1P U119 ( .A(TxData[26]), .B(TxData[27]), .C(TxData[27]), .D(
        TxData[26]), .Z(n89) );
  N1M1P U120 ( .A(TxData[28]), .Z(n87) );
  AOI22CDNM1P U121 ( .A(TxData[29]), .B(n87), .C(n87), .D(TxData[29]), .Z(n88)
         );
  EN3M1P U122 ( .A(n90), .B(n89), .C(n88), .Z(n105) );
  AOI22CDNM1P U123 ( .A(TxData[6]), .B(TxData[7]), .C(TxData[7]), .D(TxData[6]), .Z(n103) );
  AOI22CDNM1P U124 ( .A(TxData[0]), .B(TxData[1]), .C(TxData[1]), .D(TxData[0]), .Z(n95) );
  AOI22CDNM1P U125 ( .A(TxData[2]), .B(TxData[3]), .C(TxData[3]), .D(TxData[2]), .Z(n94) );
  N1M1P U126 ( .A(TxData[4]), .Z(n91) );
  AOI22CDNM1P U127 ( .A(TxData[5]), .B(n91), .C(n91), .D(TxData[5]), .Z(n92)
         );
  EN3M1P U128 ( .A(n95), .B(n94), .C(n92), .Z(n102) );
  AOI22CDNM1P U129 ( .A(TxData[15]), .B(TxData[16]), .C(TxData[16]), .D(
        TxData[15]), .Z(n99) );
  AOI22CDNM1P U130 ( .A(TxData[17]), .B(TxData[18]), .C(TxData[18]), .D(
        TxData[17]), .Z(n98) );
  N1M1P U131 ( .A(TxData[19]), .Z(n96) );
  AOI22CDNM1P U132 ( .A(TxData[23]), .B(n96), .C(n96), .D(TxData[23]), .Z(n97)
         );
  EN3M1P U133 ( .A(n99), .B(n98), .C(n97), .Z(n100) );
  EN3M1P U134 ( .A(TxData[22]), .B(TxData[14]), .C(n100), .Z(n101) );
  EN3M1P U135 ( .A(n103), .B(n102), .C(n101), .Z(n104) );
  EN3M1P U136 ( .A(n106), .B(n105), .C(n104), .Z(n113) );
  AOI22CDNM1P U137 ( .A(TxData[12]), .B(TxData[13]), .C(TxData[13]), .D(
        TxData[12]), .Z(n109) );
  AOI22CDNM1P U138 ( .A(TxData[8]), .B(TxData[9]), .C(TxData[9]), .D(TxData[8]), .Z(n108) );
  AOI22CDNM1P U139 ( .A(TxData[10]), .B(TxData[11]), .C(TxData[11]), .D(
        TxData[10]), .Z(n107) );
  EN3M1P U140 ( .A(n109), .B(n108), .C(n107), .Z(n110) );
  EN3M1P U141 ( .A(TxData[20]), .B(TxData[21]), .C(n110), .Z(n112) );
  ND2M1P U142 ( .A(n113), .B(n112), .Z(n111) );
  OAI211M1P U143 ( .A(n113), .B(n112), .C(n111), .D(n152), .Z(n114) );
  OAI21M1P U144 ( .A(n152), .B(n115), .C(n114), .Z(n144) );
  NR2M1P U145 ( .A(bitCount[3]), .B(n131), .Z(n121) );
  NR3M1P U146 ( .A(n130), .B(n128), .C(n124), .Z(n120) );
  OAI21M1P U147 ( .A(n120), .B(n131), .C(n153), .Z(n122) );
  NR2M1P U148 ( .A(n121), .B(n122), .Z(n119) );
  ND3M1P U149 ( .A(bitCount[3]), .B(n133), .C(n120), .Z(n118) );
  OAI22M1P U150 ( .A(n119), .B(n116), .C(n117), .D(n118), .Z(n146) );
  AOI22M1P U151 ( .A(bitCount[4]), .B(n119), .C(n118), .D(n117), .Z(n147) );
  AOI22M1P U152 ( .A(bitCount[3]), .B(n122), .C(n121), .D(n120), .Z(n123) );
  N1M1P U153 ( .A(n123), .Z(n148) );
  N1M1P U154 ( .A(n153), .Z(n139) );
  AOI21M1P U155 ( .A(n130), .B(n133), .C(n139), .Z(n129) );
  OA21M1P U156 ( .A(n131), .B(bitCount[1]), .C(n129), .Z(n126) );
  ND3M1P U157 ( .A(bitCount[0]), .B(bitCount[1]), .C(n133), .Z(n125) );
  AOI22M1P U158 ( .A(bitCount[2]), .B(n126), .C(n125), .D(n124), .Z(n149) );
  ND2M1P U159 ( .A(n133), .B(n128), .Z(n127) );
  OAI22M1P U160 ( .A(n129), .B(n128), .C(n130), .D(n127), .Z(n150) );
  AOI22M1P U161 ( .A(bitCount[0]), .B(n153), .C(n131), .D(n130), .Z(n151) );
  N1M1P U162 ( .A(n166), .Z(n141) );
  ND2M1P U163 ( .A(n142), .B(n141), .Z(n154) );
  NR2M1P U164 ( .A(n139), .B(n163), .Z(n132) );
  AOI211M1P U165 ( .A(n138), .B(n139), .C(n133), .D(n132), .Z(n156) );
  NR2M1P U166 ( .A(n161), .B(n145), .Z(n137) );
  N1M1P U167 ( .A(n157), .Z(n134) );
  OR3M1P U168 ( .A(n157), .B(n161), .C(n145), .Z(n136) );
  OAI211M1P U169 ( .A(n137), .B(n134), .C(n135), .D(n136), .Z(n158) );
  AO21CNM1P U170 ( .A(n159), .B(n136), .C(n135), .Z(n160) );
  AO211M1P U171 ( .A(n161), .B(n145), .C(Tx_Ready), .D(n137), .Z(n162) );
  ND3M1P U172 ( .A(n163), .B(n139), .C(n138), .Z(n140) );
endmodule


module CoreWithTxRx_Post ( Clk_r, Clk_s, Rst_n, Packet_From_Node_Valid, 
        Packet_From_Node, Packet_To_Node, Packet_To_Node_Valid, Core_Load_Ack, 
        E_Tx_Rx_Ready, E_Tx_Rx_Error, E_Tx_S_Data, E_Rx_S_Data, E_Rx_Rx_Ready, 
        E_Rx_Rx_Error, W_Tx_Rx_Ready, W_Tx_Rx_Error, W_Tx_S_Data, W_Rx_S_Data, 
        W_Rx_Rx_Ready, W_Rx_Rx_Error, S_Tx_Rx_Ready, S_Tx_Rx_Error, 
        S_Tx_S_Data, S_Rx_S_Data, S_Rx_Rx_Ready, S_Rx_Rx_Error, N_Tx_Rx_Ready, 
        N_Tx_Rx_Error, N_Tx_S_Data, N_Rx_S_Data, N_Rx_Rx_Ready, N_Rx_Rx_Error
 );
  input [31:0] Packet_From_Node;
  output [31:0] Packet_To_Node;
  input Clk_r, Clk_s, Rst_n, Packet_From_Node_Valid, E_Tx_Rx_Ready,
         E_Tx_Rx_Error, E_Rx_S_Data, W_Tx_Rx_Ready, W_Tx_Rx_Error, W_Rx_S_Data,
         S_Tx_Rx_Ready, S_Tx_Rx_Error, S_Rx_S_Data, N_Tx_Rx_Ready,
         N_Tx_Rx_Error, N_Rx_S_Data;
  output Packet_To_Node_Valid, Core_Load_Ack, E_Tx_S_Data, E_Rx_Rx_Ready,
         E_Rx_Rx_Error, W_Tx_S_Data, W_Rx_Rx_Ready, W_Rx_Rx_Error, S_Tx_S_Data,
         S_Rx_Rx_Ready, S_Rx_Rx_Error, N_Tx_S_Data, N_Rx_Rx_Ready,
         N_Rx_Rx_Error;
  wire   N_Tx_Ready, N_RxData_Valid, S_Tx_Ready, S_RxData_Valid, W_Tx_Ready,
         W_RxData_Valid, E_Tx_Ready, E_RxData_Valid, N_TxData_Valid,
         N_Core_Rcv_Ready, S_TxData_Valid, S_Core_Rcv_Ready, W_TxData_Valid,
         W_Core_Rcv_Ready, E_TxData_Valid, E_Core_Rcv_Ready;
  wire   [31:0] N_RxData;
  wire   [31:0] S_RxData;
  wire   [31:0] W_RxData;
  wire   [31:0] E_RxData;
  wire   [31:0] N_TxData;
  wire   [31:0] S_TxData;
  wire   [31:0] W_TxData;
  wire   [31:0] E_TxData;

  core routerCore ( .Clk_r(Clk_r), .Rst_n(Rst_n), .N_Tx_Ready(N_Tx_Ready), 
        .N_Tx_Error(1'b0), .N_RxData_Valid(N_RxData_Valid), .N_RxData(N_RxData), .S_Tx_Ready(S_Tx_Ready), .S_Tx_Error(1'b0), .S_RxData_Valid(S_RxData_Valid), 
        .S_RxData(S_RxData), .W_Tx_Ready(W_Tx_Ready), .W_Tx_Error(1'b0), 
        .W_RxData_Valid(W_RxData_Valid), .W_RxData(W_RxData), .E_Tx_Ready(
        E_Tx_Ready), .E_Tx_Error(1'b0), .E_RxData_Valid(E_RxData_Valid), 
        .E_RxData(E_RxData), .Packet_From_Node(Packet_From_Node), 
        .Packet_From_Node_Valid(Packet_From_Node_Valid), .N_TxData_Valid(
        N_TxData_Valid), .N_TxData(N_TxData), .N_Core_Rcv_Ready(
        N_Core_Rcv_Ready), .S_TxData_Valid(S_TxData_Valid), .S_TxData(S_TxData), .S_Core_Rcv_Ready(S_Core_Rcv_Ready), .W_TxData_Valid(W_TxData_Valid), 
        .W_TxData(W_TxData), .W_Core_Rcv_Ready(W_Core_Rcv_Ready), 
        .E_TxData_Valid(E_TxData_Valid), .E_TxData(E_TxData), 
        .E_Core_Rcv_Ready(E_Core_Rcv_Ready), .Core_Load_Ack(Core_Load_Ack), 
        .Packet_To_Node(Packet_To_Node), .Packet_To_Node_Valid(
        Packet_To_Node_Valid) );
  tx_0 E_tx ( .Clk_s(Clk_s), .Rst_n(Rst_n), .TxData_Valid(E_TxData_Valid), 
        .TxData(E_TxData), .Error_Ack(1'b0), .Rx_Ready(E_Tx_Rx_Ready), 
        .Rx_Error(1'b0), .Tx_Ready(E_Tx_Ready), .S_Data(E_Tx_S_Data) );
  rx_0 E_rx ( .Clk_s(Clk_s), .Rst_n(Rst_n), .Core_Rcv_Ready(E_Core_Rcv_Ready), 
        .S_Data(E_Rx_S_Data), .RxData_Valid(E_RxData_Valid), .RxData(E_RxData), 
        .Rx_Ready(E_Rx_Rx_Ready), .Rx_Error(E_Rx_Rx_Error) );
  tx_3 W_tx ( .Clk_s(Clk_s), .Rst_n(Rst_n), .TxData_Valid(W_TxData_Valid), 
        .TxData(W_TxData), .Error_Ack(1'b0), .Rx_Ready(W_Tx_Rx_Ready), 
        .Rx_Error(1'b0), .Tx_Ready(W_Tx_Ready), .S_Data(W_Tx_S_Data) );
  rx_3 W_rx ( .Clk_s(Clk_s), .Rst_n(Rst_n), .Core_Rcv_Ready(W_Core_Rcv_Ready), 
        .S_Data(W_Rx_S_Data), .RxData_Valid(W_RxData_Valid), .RxData(W_RxData), 
        .Rx_Ready(W_Rx_Rx_Ready), .Rx_Error(W_Rx_Rx_Error) );
  tx_2 S_tx ( .Clk_s(Clk_s), .Rst_n(Rst_n), .TxData_Valid(S_TxData_Valid), 
        .TxData(S_TxData), .Error_Ack(1'b0), .Rx_Ready(S_Tx_Rx_Ready), 
        .Rx_Error(1'b0), .Tx_Ready(S_Tx_Ready), .S_Data(S_Tx_S_Data) );
  rx_2 S_rx ( .Clk_s(Clk_s), .Rst_n(Rst_n), .Core_Rcv_Ready(S_Core_Rcv_Ready), 
        .S_Data(S_Rx_S_Data), .RxData_Valid(S_RxData_Valid), .RxData(S_RxData), 
        .Rx_Ready(S_Rx_Rx_Ready), .Rx_Error(S_Rx_Rx_Error) );
  tx_1 N_tx ( .Clk_s(Clk_s), .Rst_n(Rst_n), .TxData_Valid(N_TxData_Valid), 
        .TxData(N_TxData), .Error_Ack(1'b0), .Rx_Ready(N_Tx_Rx_Ready), 
        .Rx_Error(1'b0), .Tx_Ready(N_Tx_Ready), .S_Data(N_Tx_S_Data) );
  rx_1 N_rx ( .Clk_s(Clk_s), .Rst_n(Rst_n), .Core_Rcv_Ready(N_Core_Rcv_Ready), 
        .S_Data(N_Rx_S_Data), .RxData_Valid(N_RxData_Valid), .RxData(N_RxData), 
        .Rx_Ready(N_Rx_Rx_Ready), .Rx_Error(N_Rx_Rx_Error) );
endmodule

