library verilog;
use verilog.vl_types.all;
entity decoder_3_to_8_tb is
end decoder_3_to_8_tb;
