module cds_alias(out,in);

input in;
output out;


assign in = out;


endmodule
