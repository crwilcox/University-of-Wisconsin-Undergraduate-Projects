library verilog;
use verilog.vl_types.all;
entity p2b_adder is
end p2b_adder;
