library verilog;
use verilog.vl_types.all;
entity modulo_6_tb is
end modulo_6_tb;
