library verilog;
use verilog.vl_types.all;
entity tx_tb is
end tx_tb;
