
module Routing_State_Machine_synth ( Clk_r, Rst_n, Router_Address, Link_Config, 
        Packet_From_Link_N, Packet_From_Link_S, Packet_From_Link_W, 
        Packet_From_Link_E, Packet_From_Node, RxQueue_Empty_N, RxQueue_Empty_S, 
        RxQueue_Empty_W, RxQueue_Empty_E, TxQueue_Full_N, TxQueue_Full_S, 
        TxQueue_Full_W, TxQueue_Full_E, To_Node_Full, Node_Queue_Empty, 
        Packet_To_Link_N, Packet_To_Link_S, Packet_To_Link_W, Packet_To_Link_E, 
        Packet_To_Node, TxQueue_Write_N, TxQueue_Write_S, TxQueue_Write_W, 
        TxQueue_Write_E, To_Node_Write, RxQueue_Read_N, RxQueue_Read_S, 
        RxQueue_Read_W, RxQueue_Read_E, Node_Read );
  input [7:0] Router_Address;
  input [3:0] Link_Config;
  input [31:0] Packet_From_Link_N;
  input [31:0] Packet_From_Link_S;
  input [31:0] Packet_From_Link_W;
  input [31:0] Packet_From_Link_E;
  input [31:0] Packet_From_Node;
  output [31:0] Packet_To_Link_N;
  output [31:0] Packet_To_Link_S;
  output [31:0] Packet_To_Link_W;
  output [31:0] Packet_To_Link_E;
  output [31:0] Packet_To_Node;
  input Clk_r, Rst_n, RxQueue_Empty_N, RxQueue_Empty_S, RxQueue_Empty_W,
         RxQueue_Empty_E, TxQueue_Full_N, TxQueue_Full_S, TxQueue_Full_W,
         TxQueue_Full_E, To_Node_Full, Node_Queue_Empty;
  output TxQueue_Write_N, TxQueue_Write_S, TxQueue_Write_W, TxQueue_Write_E,
         To_Node_Write, RxQueue_Read_N, RxQueue_Read_S, RxQueue_Read_W,
         RxQueue_Read_E, Node_Read;
  wire   Packet_From_Node_31, Packet_From_Node_30, Packet_From_Node_29,
         Packet_From_Node_28, Packet_From_Node_27, Packet_From_Node_26,
         Packet_From_Node_25, Packet_From_Node_24, N44, N109, N110, N111, N112,
         N113, N114, N115, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n37, n38, n39, n40, n42, n43,
         n44, n45, n57, n107, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, \add_x_80_3/carry[7] , \add_x_80_3/carry[6] ,
         \add_x_80_3/carry[5] , \add_x_80_3/carry[4] , \add_x_80_3/carry[3] ,
         \add_x_80_3/carry[2] , n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531;
  wire   [31:0] chosenPacket;
  wire   [2:0] dataLocation;
  assign Packet_From_Node_31 = Packet_From_Node[31];
  assign Packet_From_Node_30 = Packet_From_Node[30];
  assign Packet_From_Node_29 = Packet_From_Node[29];
  assign Packet_From_Node_28 = Packet_From_Node[28];
  assign Packet_From_Node_27 = Packet_From_Node[27];
  assign Packet_From_Node_26 = Packet_From_Node[26];
  assign Packet_From_Node_25 = Packet_From_Node[25];
  assign Packet_From_Node_24 = Packet_From_Node[24];

  FD4QM1P \Packet_To_Node_reg[16]  ( .D(n25), .CP(Clk_r), .SD(Rst_n), .Q(
        Packet_To_Node[16]) );
  FD4QM1P \Packet_To_Node_reg[17]  ( .D(n26), .CP(Clk_r), .SD(Rst_n), .Q(
        Packet_To_Node[17]) );
  FD4QM1P \Packet_To_Node_reg[18]  ( .D(n27), .CP(Clk_r), .SD(Rst_n), .Q(
        Packet_To_Node[18]) );
  FD4QM1P \Packet_To_Node_reg[19]  ( .D(n28), .CP(Clk_r), .SD(Rst_n), .Q(
        Packet_To_Node[19]) );
  FD4QM1P \Packet_To_Node_reg[20]  ( .D(n29), .CP(Clk_r), .SD(Rst_n), .Q(
        Packet_To_Node[20]) );
  FD4QM1P \Packet_To_Node_reg[21]  ( .D(n30), .CP(Clk_r), .SD(Rst_n), .Q(
        Packet_To_Node[21]) );
  FD4QM1P \Packet_To_Node_reg[22]  ( .D(n31), .CP(Clk_r), .SD(Rst_n), .Q(
        Packet_To_Node[22]) );
  FD4QM1P \Packet_To_Node_reg[23]  ( .D(n32), .CP(Clk_r), .SD(Rst_n), .Q(
        Packet_To_Node[23]) );
  FD2QM1P To_Node_Write_reg ( .D(n261), .CP(Clk_r), .CD(Rst_n), .Q(
        To_Node_Write) );
  FD2LQM1P \Packet_To_Node_reg[31]  ( .D(n491), .LD(n327), .CP(Clk_r), .CD(
        Rst_n), .Q(n5) );
  FD2LQM1P \Packet_To_Node_reg[30]  ( .D(n42), .LD(n327), .CP(Clk_r), .CD(
        Rst_n), .Q(n4) );
  FD2LQM1P \Packet_To_Node_reg[29]  ( .D(n43), .LD(n328), .CP(Clk_r), .CD(
        Rst_n), .Q(n3) );
  FD2LQM1P \Packet_To_Node_reg[27]  ( .D(n44), .LD(n327), .CP(Clk_r), .CD(
        Rst_n), .Q(n2) );
  FD4QM1P \Packet_To_Node_reg[26]  ( .D(n34), .CP(Clk_r), .SD(Rst_n), .Q(
        Packet_To_Node[26]) );
  FD2LQM1P \Packet_To_Node_reg[25]  ( .D(n45), .LD(n327), .CP(Clk_r), .CD(
        Rst_n), .Q(n1) );
  FD1LQM1P \Packet_To_Link_N_reg[31]  ( .D(chosenPacket[31]), .LD(n333), .CP(
        Clk_r), .Q(Packet_To_Link_N[31]) );
  FD1LQM1P \Packet_To_Link_N_reg[30]  ( .D(chosenPacket[30]), .LD(n333), .CP(
        Clk_r), .Q(Packet_To_Link_N[30]) );
  FD1LQM1P \Packet_To_Link_N_reg[29]  ( .D(chosenPacket[29]), .LD(n333), .CP(
        Clk_r), .Q(Packet_To_Link_N[29]) );
  FD1LQM1P \Packet_To_Link_N_reg[27]  ( .D(chosenPacket[27]), .LD(n333), .CP(
        Clk_r), .Q(Packet_To_Link_N[27]) );
  FD1LQM1P \Packet_To_Link_N_reg[25]  ( .D(chosenPacket[25]), .LD(n333), .CP(
        Clk_r), .Q(Packet_To_Link_N[25]) );
  FD1LQM1P \Packet_To_Link_N_reg[16]  ( .D(n310), .LD(n333), .CP(Clk_r), .Q(
        Packet_To_Link_N[16]) );
  FD1LQM1P \Packet_To_Link_N_reg[17]  ( .D(N109), .LD(n333), .CP(Clk_r), .Q(
        Packet_To_Link_N[17]) );
  FD1LQM1P \Packet_To_Link_N_reg[18]  ( .D(N110), .LD(n333), .CP(Clk_r), .Q(
        Packet_To_Link_N[18]) );
  FD1LQM1P \Packet_To_Link_N_reg[19]  ( .D(N111), .LD(n333), .CP(Clk_r), .Q(
        Packet_To_Link_N[19]) );
  FD1LQM1P \Packet_To_Link_N_reg[20]  ( .D(N112), .LD(n333), .CP(Clk_r), .Q(
        Packet_To_Link_N[20]) );
  FD1LQM1P \Packet_To_Link_N_reg[21]  ( .D(N113), .LD(n333), .CP(Clk_r), .Q(
        Packet_To_Link_N[21]) );
  FD1LQM1P \Packet_To_Link_N_reg[22]  ( .D(N114), .LD(n333), .CP(Clk_r), .Q(
        Packet_To_Link_N[22]) );
  FD1LQM1P \Packet_To_Link_N_reg[23]  ( .D(N115), .LD(n333), .CP(Clk_r), .Q(
        Packet_To_Link_N[23]) );
  FD1LQM1P \Packet_To_Link_N_reg[26]  ( .D(chosenPacket[26]), .LD(n333), .CP(
        Clk_r), .Q(Packet_To_Link_N[26]) );
  FD1LQM1P \Packet_To_Link_N_reg[28]  ( .D(chosenPacket[28]), .LD(n333), .CP(
        Clk_r), .Q(Packet_To_Link_N[28]) );
  FD1LQM1P \Packet_To_Link_S_reg[31]  ( .D(chosenPacket[31]), .LD(n330), .CP(
        Clk_r), .Q(Packet_To_Link_S[31]) );
  FD1LQM1P \Packet_To_Link_S_reg[30]  ( .D(chosenPacket[30]), .LD(n330), .CP(
        Clk_r), .Q(Packet_To_Link_S[30]) );
  FD1LQM1P \Packet_To_Link_S_reg[29]  ( .D(chosenPacket[29]), .LD(n330), .CP(
        Clk_r), .Q(Packet_To_Link_S[29]) );
  FD1LQM1P \Packet_To_Link_S_reg[27]  ( .D(chosenPacket[27]), .LD(n330), .CP(
        Clk_r), .Q(Packet_To_Link_S[27]) );
  FD1LQM1P \Packet_To_Link_S_reg[25]  ( .D(chosenPacket[25]), .LD(n330), .CP(
        Clk_r), .Q(Packet_To_Link_S[25]) );
  FD1LQM1P \Packet_To_Link_S_reg[16]  ( .D(n310), .LD(n330), .CP(Clk_r), .Q(
        Packet_To_Link_S[16]) );
  FD1LQM1P \Packet_To_Link_S_reg[17]  ( .D(N109), .LD(n330), .CP(Clk_r), .Q(
        Packet_To_Link_S[17]) );
  FD1LQM1P \Packet_To_Link_S_reg[18]  ( .D(N110), .LD(n330), .CP(Clk_r), .Q(
        Packet_To_Link_S[18]) );
  FD1LQM1P \Packet_To_Link_S_reg[19]  ( .D(N111), .LD(n330), .CP(Clk_r), .Q(
        Packet_To_Link_S[19]) );
  FD1LQM1P \Packet_To_Link_S_reg[20]  ( .D(N112), .LD(n330), .CP(Clk_r), .Q(
        Packet_To_Link_S[20]) );
  FD1LQM1P \Packet_To_Link_S_reg[21]  ( .D(N113), .LD(n331), .CP(Clk_r), .Q(
        Packet_To_Link_S[21]) );
  FD1LQM1P \Packet_To_Link_S_reg[22]  ( .D(N114), .LD(n331), .CP(Clk_r), .Q(
        Packet_To_Link_S[22]) );
  FD1LQM1P \Packet_To_Link_S_reg[23]  ( .D(n303), .LD(n331), .CP(Clk_r), .Q(
        Packet_To_Link_S[23]) );
  FD1LQM1P \Packet_To_Link_S_reg[26]  ( .D(chosenPacket[26]), .LD(n331), .CP(
        Clk_r), .Q(Packet_To_Link_S[26]) );
  FD1LQM1P \Packet_To_Link_S_reg[28]  ( .D(chosenPacket[28]), .LD(n331), .CP(
        Clk_r), .Q(Packet_To_Link_S[28]) );
  FD1LQM1P \Packet_To_Link_W_reg[31]  ( .D(chosenPacket[31]), .LD(n312), .CP(
        Clk_r), .Q(Packet_To_Link_W[31]) );
  FD1LQM1P \Packet_To_Link_W_reg[30]  ( .D(chosenPacket[30]), .LD(n302), .CP(
        Clk_r), .Q(Packet_To_Link_W[30]) );
  FD1LQM1P \Packet_To_Link_W_reg[29]  ( .D(chosenPacket[29]), .LD(n302), .CP(
        Clk_r), .Q(Packet_To_Link_W[29]) );
  FD1LQM1P \Packet_To_Link_W_reg[27]  ( .D(chosenPacket[27]), .LD(n313), .CP(
        Clk_r), .Q(Packet_To_Link_W[27]) );
  FD1LQM1P \Packet_To_Link_W_reg[25]  ( .D(chosenPacket[25]), .LD(n312), .CP(
        Clk_r), .Q(Packet_To_Link_W[25]) );
  FD1LQM1P \Packet_To_Link_W_reg[16]  ( .D(n310), .LD(n313), .CP(Clk_r), .Q(
        Packet_To_Link_W[16]) );
  FD1LQM1P \Packet_To_Link_W_reg[17]  ( .D(N109), .LD(n312), .CP(Clk_r), .Q(
        Packet_To_Link_W[17]) );
  FD1LQM1P \Packet_To_Link_W_reg[18]  ( .D(N110), .LD(n313), .CP(Clk_r), .Q(
        Packet_To_Link_W[18]) );
  FD1LQM1P \Packet_To_Link_W_reg[19]  ( .D(N111), .LD(n312), .CP(Clk_r), .Q(
        Packet_To_Link_W[19]) );
  FD1LQM1P \Packet_To_Link_W_reg[20]  ( .D(N112), .LD(n313), .CP(Clk_r), .Q(
        Packet_To_Link_W[20]) );
  FD1LQM1P \Packet_To_Link_W_reg[21]  ( .D(N113), .LD(n302), .CP(Clk_r), .Q(
        Packet_To_Link_W[21]) );
  FD1LQM1P \Packet_To_Link_W_reg[22]  ( .D(N114), .LD(n313), .CP(Clk_r), .Q(
        Packet_To_Link_W[22]) );
  FD1LQM1P \Packet_To_Link_W_reg[23]  ( .D(n303), .LD(n302), .CP(Clk_r), .Q(
        Packet_To_Link_W[23]) );
  FD1LQM1P \Packet_To_Link_W_reg[26]  ( .D(chosenPacket[26]), .LD(n302), .CP(
        Clk_r), .Q(Packet_To_Link_W[26]) );
  FD1LQM1P \Packet_To_Link_W_reg[28]  ( .D(chosenPacket[28]), .LD(n302), .CP(
        Clk_r), .Q(Packet_To_Link_W[28]) );
  FD1LQM1P \Packet_To_Link_E_reg[31]  ( .D(chosenPacket[31]), .LD(n316), .CP(
        Clk_r), .Q(Packet_To_Link_E[31]) );
  FD1LQM1P \Packet_To_Link_E_reg[30]  ( .D(chosenPacket[30]), .LD(n315), .CP(
        Clk_r), .Q(Packet_To_Link_E[30]) );
  FD1LQM1P \Packet_To_Link_E_reg[29]  ( .D(chosenPacket[29]), .LD(n316), .CP(
        Clk_r), .Q(Packet_To_Link_E[29]) );
  FD1LQM1P \Packet_To_Link_E_reg[27]  ( .D(chosenPacket[27]), .LD(n317), .CP(
        Clk_r), .Q(Packet_To_Link_E[27]) );
  FD1LQM1P \Packet_To_Link_E_reg[25]  ( .D(chosenPacket[25]), .LD(n316), .CP(
        Clk_r), .Q(Packet_To_Link_E[25]) );
  FD1LQM1P \Packet_To_Link_E_reg[16]  ( .D(n310), .LD(n315), .CP(Clk_r), .Q(
        Packet_To_Link_E[16]) );
  FD1LQM1P \Packet_To_Link_E_reg[17]  ( .D(N109), .LD(n315), .CP(Clk_r), .Q(
        Packet_To_Link_E[17]) );
  FD1LQM1P \Packet_To_Link_E_reg[18]  ( .D(N110), .LD(n317), .CP(Clk_r), .Q(
        Packet_To_Link_E[18]) );
  FD1LQM1P \Packet_To_Link_E_reg[19]  ( .D(N111), .LD(n317), .CP(Clk_r), .Q(
        Packet_To_Link_E[19]) );
  FD1LQM1P \Packet_To_Link_E_reg[20]  ( .D(N112), .LD(n316), .CP(Clk_r), .Q(
        Packet_To_Link_E[20]) );
  FD1LQM1P \Packet_To_Link_E_reg[21]  ( .D(N113), .LD(n317), .CP(Clk_r), .Q(
        Packet_To_Link_E[21]) );
  FD1LQM1P \Packet_To_Link_E_reg[22]  ( .D(N114), .LD(n316), .CP(Clk_r), .Q(
        Packet_To_Link_E[22]) );
  FD1LQM1P \Packet_To_Link_E_reg[23]  ( .D(n303), .LD(n315), .CP(Clk_r), .Q(
        Packet_To_Link_E[23]) );
  FD1LQM1P \Packet_To_Link_E_reg[26]  ( .D(chosenPacket[26]), .LD(n316), .CP(
        Clk_r), .Q(Packet_To_Link_E[26]) );
  FD1LQM1P \Packet_To_Link_E_reg[28]  ( .D(chosenPacket[28]), .LD(n317), .CP(
        Clk_r), .Q(Packet_To_Link_E[28]) );
  FD1LQM1P \Packet_To_Link_E_reg[24]  ( .D(chosenPacket[24]), .LD(n316), .CP(
        Clk_r), .Q(Packet_To_Link_E[24]) );
  FD4QM1P \Packet_To_Node_reg[24]  ( .D(n33), .CP(Clk_r), .SD(Rst_n), .Q(
        Packet_To_Node[24]) );
  FD1LQM1P \Packet_To_Link_W_reg[24]  ( .D(chosenPacket[24]), .LD(n312), .CP(
        Clk_r), .Q(Packet_To_Link_W[24]) );
  FD1LQM1P \Packet_To_Link_N_reg[24]  ( .D(chosenPacket[24]), .LD(n333), .CP(
        Clk_r), .Q(Packet_To_Link_N[24]) );
  FD1LQM1P \Packet_To_Link_S_reg[24]  ( .D(chosenPacket[24]), .LD(n331), .CP(
        Clk_r), .Q(Packet_To_Link_S[24]) );
  FD1QM1P \chosenPacket_reg[15]  ( .D(n271), .CP(Clk_r), .Q(chosenPacket[15])
         );
  FD1LQM1P \Packet_To_Link_E_reg[15]  ( .D(chosenPacket[15]), .LD(n315), .CP(
        Clk_r), .Q(Packet_To_Link_E[15]) );
  FD4QM1P \Packet_To_Node_reg[15]  ( .D(n24), .CP(Clk_r), .SD(Rst_n), .Q(
        Packet_To_Node[15]) );
  FD1LQM1P \Packet_To_Link_W_reg[15]  ( .D(chosenPacket[15]), .LD(n312), .CP(
        Clk_r), .Q(Packet_To_Link_W[15]) );
  FD1LQM1P \Packet_To_Link_N_reg[15]  ( .D(chosenPacket[15]), .LD(n333), .CP(
        Clk_r), .Q(Packet_To_Link_N[15]) );
  FD1LQM1P \Packet_To_Link_S_reg[15]  ( .D(chosenPacket[15]), .LD(n331), .CP(
        Clk_r), .Q(Packet_To_Link_S[15]) );
  FD1QM1P \chosenPacket_reg[14]  ( .D(n272), .CP(Clk_r), .Q(chosenPacket[14])
         );
  FD1LQM1P \Packet_To_Link_E_reg[14]  ( .D(chosenPacket[14]), .LD(n315), .CP(
        Clk_r), .Q(Packet_To_Link_E[14]) );
  FD4QM1P \Packet_To_Node_reg[14]  ( .D(n23), .CP(Clk_r), .SD(Rst_n), .Q(
        Packet_To_Node[14]) );
  FD1LQM1P \Packet_To_Link_W_reg[14]  ( .D(chosenPacket[14]), .LD(n302), .CP(
        Clk_r), .Q(Packet_To_Link_W[14]) );
  FD1LQM1P \Packet_To_Link_N_reg[14]  ( .D(chosenPacket[14]), .LD(n333), .CP(
        Clk_r), .Q(Packet_To_Link_N[14]) );
  FD1LQM1P \Packet_To_Link_S_reg[14]  ( .D(chosenPacket[14]), .LD(n331), .CP(
        Clk_r), .Q(Packet_To_Link_S[14]) );
  FD1QM1P \chosenPacket_reg[13]  ( .D(n273), .CP(Clk_r), .Q(chosenPacket[13])
         );
  FD1LQM1P \Packet_To_Link_E_reg[13]  ( .D(chosenPacket[13]), .LD(n317), .CP(
        Clk_r), .Q(Packet_To_Link_E[13]) );
  FD4QM1P \Packet_To_Node_reg[13]  ( .D(n22), .CP(Clk_r), .SD(Rst_n), .Q(
        Packet_To_Node[13]) );
  FD1LQM1P \Packet_To_Link_W_reg[13]  ( .D(chosenPacket[13]), .LD(n313), .CP(
        Clk_r), .Q(Packet_To_Link_W[13]) );
  FD1LQM1P \Packet_To_Link_N_reg[13]  ( .D(chosenPacket[13]), .LD(n333), .CP(
        Clk_r), .Q(Packet_To_Link_N[13]) );
  FD1LQM1P \Packet_To_Link_S_reg[13]  ( .D(chosenPacket[13]), .LD(n331), .CP(
        Clk_r), .Q(Packet_To_Link_S[13]) );
  FD1QM1P \chosenPacket_reg[12]  ( .D(n274), .CP(Clk_r), .Q(chosenPacket[12])
         );
  FD1LQM1P \Packet_To_Link_E_reg[12]  ( .D(chosenPacket[12]), .LD(n317), .CP(
        Clk_r), .Q(Packet_To_Link_E[12]) );
  FD4QM1P \Packet_To_Node_reg[12]  ( .D(n21), .CP(Clk_r), .SD(Rst_n), .Q(
        Packet_To_Node[12]) );
  FD1LQM1P \Packet_To_Link_W_reg[12]  ( .D(chosenPacket[12]), .LD(n312), .CP(
        Clk_r), .Q(Packet_To_Link_W[12]) );
  FD1LQM1P \Packet_To_Link_N_reg[12]  ( .D(chosenPacket[12]), .LD(n333), .CP(
        Clk_r), .Q(Packet_To_Link_N[12]) );
  FD1LQM1P \Packet_To_Link_S_reg[12]  ( .D(chosenPacket[12]), .LD(n331), .CP(
        Clk_r), .Q(Packet_To_Link_S[12]) );
  FD1QM1P \chosenPacket_reg[11]  ( .D(n275), .CP(Clk_r), .Q(chosenPacket[11])
         );
  FD1LQM1P \Packet_To_Link_E_reg[11]  ( .D(chosenPacket[11]), .LD(n315), .CP(
        Clk_r), .Q(Packet_To_Link_E[11]) );
  FD4QM1P \Packet_To_Node_reg[11]  ( .D(n20), .CP(Clk_r), .SD(Rst_n), .Q(
        Packet_To_Node[11]) );
  FD1LQM1P \Packet_To_Link_W_reg[11]  ( .D(chosenPacket[11]), .LD(n312), .CP(
        Clk_r), .Q(Packet_To_Link_W[11]) );
  FD1LQM1P \Packet_To_Link_N_reg[11]  ( .D(chosenPacket[11]), .LD(n333), .CP(
        Clk_r), .Q(Packet_To_Link_N[11]) );
  FD1LQM1P \Packet_To_Link_S_reg[11]  ( .D(chosenPacket[11]), .LD(n332), .CP(
        Clk_r), .Q(Packet_To_Link_S[11]) );
  FD1QM1P \chosenPacket_reg[10]  ( .D(n276), .CP(Clk_r), .Q(chosenPacket[10])
         );
  FD1LQM1P \Packet_To_Link_E_reg[10]  ( .D(chosenPacket[10]), .LD(n316), .CP(
        Clk_r), .Q(Packet_To_Link_E[10]) );
  FD4QM1P \Packet_To_Node_reg[10]  ( .D(n19), .CP(Clk_r), .SD(Rst_n), .Q(
        Packet_To_Node[10]) );
  FD1LQM1P \Packet_To_Link_W_reg[10]  ( .D(chosenPacket[10]), .LD(n313), .CP(
        Clk_r), .Q(Packet_To_Link_W[10]) );
  FD1LQM1P \Packet_To_Link_N_reg[10]  ( .D(chosenPacket[10]), .LD(n333), .CP(
        Clk_r), .Q(Packet_To_Link_N[10]) );
  FD1LQM1P \Packet_To_Link_S_reg[10]  ( .D(chosenPacket[10]), .LD(n332), .CP(
        Clk_r), .Q(Packet_To_Link_S[10]) );
  FD1QM1P \chosenPacket_reg[9]  ( .D(n277), .CP(Clk_r), .Q(chosenPacket[9]) );
  FD1LQM1P \Packet_To_Link_E_reg[9]  ( .D(chosenPacket[9]), .LD(n317), .CP(
        Clk_r), .Q(Packet_To_Link_E[9]) );
  FD4QM1P \Packet_To_Node_reg[9]  ( .D(n18), .CP(Clk_r), .SD(Rst_n), .Q(
        Packet_To_Node[9]) );
  FD1LQM1P \Packet_To_Link_W_reg[9]  ( .D(chosenPacket[9]), .LD(n312), .CP(
        Clk_r), .Q(Packet_To_Link_W[9]) );
  FD1LQM1P \Packet_To_Link_N_reg[9]  ( .D(chosenPacket[9]), .LD(n333), .CP(
        Clk_r), .Q(Packet_To_Link_N[9]) );
  FD1LQM1P \Packet_To_Link_S_reg[9]  ( .D(chosenPacket[9]), .LD(n332), .CP(
        Clk_r), .Q(Packet_To_Link_S[9]) );
  FD1QM1P \chosenPacket_reg[8]  ( .D(n278), .CP(Clk_r), .Q(chosenPacket[8]) );
  FD1LQM1P \Packet_To_Link_E_reg[8]  ( .D(chosenPacket[8]), .LD(n316), .CP(
        Clk_r), .Q(Packet_To_Link_E[8]) );
  FD4QM1P \Packet_To_Node_reg[8]  ( .D(n17), .CP(Clk_r), .SD(Rst_n), .Q(
        Packet_To_Node[8]) );
  FD1LQM1P \Packet_To_Link_W_reg[8]  ( .D(chosenPacket[8]), .LD(n302), .CP(
        Clk_r), .Q(Packet_To_Link_W[8]) );
  FD1LQM1P \Packet_To_Link_N_reg[8]  ( .D(chosenPacket[8]), .LD(n333), .CP(
        Clk_r), .Q(Packet_To_Link_N[8]) );
  FD1LQM1P \Packet_To_Link_S_reg[8]  ( .D(chosenPacket[8]), .LD(n332), .CP(
        Clk_r), .Q(Packet_To_Link_S[8]) );
  FD1QM1P \chosenPacket_reg[7]  ( .D(n279), .CP(Clk_r), .Q(chosenPacket[7]) );
  FD1LQM1P \Packet_To_Link_E_reg[7]  ( .D(chosenPacket[7]), .LD(n315), .CP(
        Clk_r), .Q(Packet_To_Link_E[7]) );
  FD4QM1P \Packet_To_Node_reg[7]  ( .D(n16), .CP(Clk_r), .SD(Rst_n), .Q(
        Packet_To_Node[7]) );
  FD1LQM1P \Packet_To_Link_W_reg[7]  ( .D(chosenPacket[7]), .LD(n313), .CP(
        Clk_r), .Q(Packet_To_Link_W[7]) );
  FD1LQM1P \Packet_To_Link_N_reg[7]  ( .D(chosenPacket[7]), .LD(n333), .CP(
        Clk_r), .Q(Packet_To_Link_N[7]) );
  FD1LQM1P \Packet_To_Link_S_reg[7]  ( .D(chosenPacket[7]), .LD(n332), .CP(
        Clk_r), .Q(Packet_To_Link_S[7]) );
  FD1QM1P \chosenPacket_reg[6]  ( .D(n280), .CP(Clk_r), .Q(chosenPacket[6]) );
  FD1LQM1P \Packet_To_Link_E_reg[6]  ( .D(chosenPacket[6]), .LD(n315), .CP(
        Clk_r), .Q(Packet_To_Link_E[6]) );
  FD4QM1P \Packet_To_Node_reg[6]  ( .D(n15), .CP(Clk_r), .SD(Rst_n), .Q(
        Packet_To_Node[6]) );
  FD1LQM1P \Packet_To_Link_W_reg[6]  ( .D(chosenPacket[6]), .LD(n313), .CP(
        Clk_r), .Q(Packet_To_Link_W[6]) );
  FD1LQM1P \Packet_To_Link_N_reg[6]  ( .D(chosenPacket[6]), .LD(n333), .CP(
        Clk_r), .Q(Packet_To_Link_N[6]) );
  FD1LQM1P \Packet_To_Link_S_reg[6]  ( .D(chosenPacket[6]), .LD(n332), .CP(
        Clk_r), .Q(Packet_To_Link_S[6]) );
  FD1QM1P \chosenPacket_reg[5]  ( .D(n281), .CP(Clk_r), .Q(chosenPacket[5]) );
  FD1LQM1P \Packet_To_Link_E_reg[5]  ( .D(chosenPacket[5]), .LD(n317), .CP(
        Clk_r), .Q(Packet_To_Link_E[5]) );
  FD4QM1P \Packet_To_Node_reg[5]  ( .D(n14), .CP(Clk_r), .SD(Rst_n), .Q(
        Packet_To_Node[5]) );
  FD1LQM1P \Packet_To_Link_W_reg[5]  ( .D(chosenPacket[5]), .LD(n302), .CP(
        Clk_r), .Q(Packet_To_Link_W[5]) );
  FD1LQM1P \Packet_To_Link_N_reg[5]  ( .D(chosenPacket[5]), .LD(n333), .CP(
        Clk_r), .Q(Packet_To_Link_N[5]) );
  FD1LQM1P \Packet_To_Link_S_reg[5]  ( .D(chosenPacket[5]), .LD(n332), .CP(
        Clk_r), .Q(Packet_To_Link_S[5]) );
  FD1QM1P \chosenPacket_reg[4]  ( .D(n282), .CP(Clk_r), .Q(chosenPacket[4]) );
  FD1LQM1P \Packet_To_Link_E_reg[4]  ( .D(chosenPacket[4]), .LD(n317), .CP(
        Clk_r), .Q(Packet_To_Link_E[4]) );
  FD4QM1P \Packet_To_Node_reg[4]  ( .D(n13), .CP(Clk_r), .SD(Rst_n), .Q(
        Packet_To_Node[4]) );
  FD1LQM1P \Packet_To_Link_W_reg[4]  ( .D(chosenPacket[4]), .LD(n313), .CP(
        Clk_r), .Q(Packet_To_Link_W[4]) );
  FD1LQM1P \Packet_To_Link_N_reg[4]  ( .D(chosenPacket[4]), .LD(n333), .CP(
        Clk_r), .Q(Packet_To_Link_N[4]) );
  FD1LQM1P \Packet_To_Link_S_reg[4]  ( .D(chosenPacket[4]), .LD(n332), .CP(
        Clk_r), .Q(Packet_To_Link_S[4]) );
  FD1QM1P \chosenPacket_reg[3]  ( .D(n283), .CP(Clk_r), .Q(chosenPacket[3]) );
  FD1LQM1P \Packet_To_Link_E_reg[3]  ( .D(chosenPacket[3]), .LD(n316), .CP(
        Clk_r), .Q(Packet_To_Link_E[3]) );
  FD4QM1P \Packet_To_Node_reg[3]  ( .D(n12), .CP(Clk_r), .SD(Rst_n), .Q(
        Packet_To_Node[3]) );
  FD1LQM1P \Packet_To_Link_W_reg[3]  ( .D(chosenPacket[3]), .LD(n312), .CP(
        Clk_r), .Q(Packet_To_Link_W[3]) );
  FD1LQM1P \Packet_To_Link_N_reg[3]  ( .D(chosenPacket[3]), .LD(n333), .CP(
        Clk_r), .Q(Packet_To_Link_N[3]) );
  FD1LQM1P \Packet_To_Link_S_reg[3]  ( .D(chosenPacket[3]), .LD(n332), .CP(
        Clk_r), .Q(Packet_To_Link_S[3]) );
  FD1QM1P \chosenPacket_reg[2]  ( .D(n284), .CP(Clk_r), .Q(chosenPacket[2]) );
  FD1LQM1P \Packet_To_Link_E_reg[2]  ( .D(chosenPacket[2]), .LD(n315), .CP(
        Clk_r), .Q(Packet_To_Link_E[2]) );
  FD4QM1P \Packet_To_Node_reg[2]  ( .D(n11), .CP(Clk_r), .SD(Rst_n), .Q(
        Packet_To_Node[2]) );
  FD1LQM1P \Packet_To_Link_W_reg[2]  ( .D(chosenPacket[2]), .LD(n302), .CP(
        Clk_r), .Q(Packet_To_Link_W[2]) );
  FD1LQM1P \Packet_To_Link_N_reg[2]  ( .D(chosenPacket[2]), .LD(n333), .CP(
        Clk_r), .Q(Packet_To_Link_N[2]) );
  FD1LQM1P \Packet_To_Link_S_reg[2]  ( .D(chosenPacket[2]), .LD(n332), .CP(
        Clk_r), .Q(Packet_To_Link_S[2]) );
  FD1QM1P \chosenPacket_reg[1]  ( .D(n285), .CP(Clk_r), .Q(chosenPacket[1]) );
  FD1LQM1P \Packet_To_Link_E_reg[1]  ( .D(chosenPacket[1]), .LD(n316), .CP(
        Clk_r), .Q(Packet_To_Link_E[1]) );
  FD4QM1P \Packet_To_Node_reg[1]  ( .D(n10), .CP(Clk_r), .SD(Rst_n), .Q(
        Packet_To_Node[1]) );
  FD1LQM1P \Packet_To_Link_W_reg[1]  ( .D(chosenPacket[1]), .LD(n312), .CP(
        Clk_r), .Q(Packet_To_Link_W[1]) );
  FD1LQM1P \Packet_To_Link_N_reg[1]  ( .D(chosenPacket[1]), .LD(n333), .CP(
        Clk_r), .Q(Packet_To_Link_N[1]) );
  FD1LQM1P \Packet_To_Link_S_reg[1]  ( .D(chosenPacket[1]), .LD(n331), .CP(
        Clk_r), .Q(Packet_To_Link_S[1]) );
  FD1QM1P \chosenPacket_reg[0]  ( .D(n286), .CP(Clk_r), .Q(chosenPacket[0]) );
  FD1LQM1P \Packet_To_Link_E_reg[0]  ( .D(chosenPacket[0]), .LD(n316), .CP(
        Clk_r), .Q(Packet_To_Link_E[0]) );
  FD4QM1P \Packet_To_Node_reg[0]  ( .D(n9), .CP(Clk_r), .SD(Rst_n), .Q(
        Packet_To_Node[0]) );
  FD1LQM1P \Packet_To_Link_W_reg[0]  ( .D(chosenPacket[0]), .LD(n313), .CP(
        Clk_r), .Q(Packet_To_Link_W[0]) );
  FD1LQM1P \Packet_To_Link_N_reg[0]  ( .D(chosenPacket[0]), .LD(n333), .CP(
        Clk_r), .Q(Packet_To_Link_N[0]) );
  FD1LQM1P \Packet_To_Link_S_reg[0]  ( .D(chosenPacket[0]), .LD(n330), .CP(
        Clk_r), .Q(Packet_To_Link_S[0]) );
  FD1QM1P \chosenPacket_reg[23]  ( .D(n262), .CP(Clk_r), .Q(chosenPacket[23])
         );
  FD1QM1P \chosenPacket_reg[18]  ( .D(n258), .CP(Clk_r), .Q(chosenPacket[18])
         );
  FD1QM1P \chosenPacket_reg[19]  ( .D(n257), .CP(Clk_r), .Q(chosenPacket[19])
         );
  FD1QM1P \chosenPacket_reg[20]  ( .D(n256), .CP(Clk_r), .Q(chosenPacket[20])
         );
  FD1QM1P \chosenPacket_reg[21]  ( .D(n255), .CP(Clk_r), .Q(chosenPacket[21])
         );
  FD1QM1P \chosenPacket_reg[22]  ( .D(n254), .CP(Clk_r), .Q(chosenPacket[22])
         );
  FD2QM1P \TxQueue_Write_reg[3]  ( .D(n253), .CP(Clk_r), .CD(Rst_n), .Q(
        TxQueue_Write_N) );
  FD2QM1P \TxQueue_Write_reg[2]  ( .D(n252), .CP(Clk_r), .CD(Rst_n), .Q(
        TxQueue_Write_S) );
  FD2QM1P \TxQueue_Write_reg[1]  ( .D(n251), .CP(Clk_r), .CD(Rst_n), .Q(
        TxQueue_Write_W) );
  FD2QM1P \TxQueue_Write_reg[0]  ( .D(n250), .CP(Clk_r), .CD(Rst_n), .Q(
        TxQueue_Write_E) );
  FD2QM1P \RxQueue_Read_reg[4]  ( .D(n245), .CP(Clk_r), .CD(Rst_n), .Q(
        Node_Read) );
  FD2QM1P \RxQueue_Read_reg[3]  ( .D(n246), .CP(Clk_r), .CD(Rst_n), .Q(
        RxQueue_Read_N) );
  FD2QM1P \RxQueue_Read_reg[2]  ( .D(n247), .CP(Clk_r), .CD(Rst_n), .Q(
        RxQueue_Read_S) );
  FD2QM1P \RxQueue_Read_reg[1]  ( .D(n248), .CP(Clk_r), .CD(Rst_n), .Q(
        RxQueue_Read_W) );
  FD2QM1P \RxQueue_Read_reg[0]  ( .D(n249), .CP(Clk_r), .CD(Rst_n), .Q(
        RxQueue_Read_E) );
  FD2LQM3P \dataLocation_reg[2]  ( .D(n57), .LD(n8), .CP(Clk_r), .CD(Rst_n), 
        .Q(n6) );
  FD1QM1P \chosenPacket_reg[28]  ( .D(n266), .CP(Clk_r), .Q(chosenPacket[28])
         );
  FD1QM1P \chosenPacket_reg[26]  ( .D(n268), .CP(Clk_r), .Q(chosenPacket[26])
         );
  FD1QM3P \chosenPacket_reg[29]  ( .D(n265), .CP(Clk_r), .Q(chosenPacket[29])
         );
  FD1QM1P \chosenPacket_reg[30]  ( .D(n264), .CP(Clk_r), .Q(chosenPacket[30])
         );
  FD1QM3P \chosenPacket_reg[25]  ( .D(n269), .CP(Clk_r), .Q(chosenPacket[25])
         );
  FD1QM3P \chosenPacket_reg[24]  ( .D(n270), .CP(Clk_r), .Q(chosenPacket[24])
         );
  FD1QM1P \chosenPacket_reg[31]  ( .D(n263), .CP(Clk_r), .Q(chosenPacket[31])
         );
  FD4QM1P \nextStage_reg[0]  ( .D(n7), .CP(Clk_r), .SD(Rst_n), .Q(n8) );
  FD1QM3P \chosenPacket_reg[17]  ( .D(n259), .CP(Clk_r), .Q(chosenPacket[17])
         );
  FD2LQM3P \dataLocation_reg[1]  ( .D(N44), .LD(n8), .CP(Clk_r), .CD(Rst_n), 
        .Q(dataLocation[1]) );
  FD2LQM1P \dataLocation_reg[0]  ( .D(n488), .LD(n8), .CP(Clk_r), .CD(Rst_n), 
        .Q(dataLocation[0]) );
  FD2LQM1P \Packet_To_Node_reg[28]  ( .D(n514), .LD(n107), .CP(Clk_r), .CD(
        Rst_n), .Q(n304) );
  FD1QM3P \chosenPacket_reg[27]  ( .D(n267), .CP(Clk_r), .Q(chosenPacket[27])
         );
  FD1QM8P \chosenPacket_reg[16]  ( .D(n260), .CP(Clk_r), .Q(chosenPacket[16])
         );
  NR2M2P U294 ( .A(n477), .B(n377), .Z(n474) );
  AND2M2P U295 ( .A(n6), .B(dataLocation[0]), .Z(n340) );
  BUFM2P U296 ( .A(n478), .Z(n324) );
  BUFM2P U297 ( .A(n478), .Z(n325) );
  BUFM6P U298 ( .A(n476), .Z(n306) );
  BUFM2P U299 ( .A(n478), .Z(n326) );
  BUFM4P U300 ( .A(n473), .Z(n305) );
  N1M1P U301 ( .A(chosenPacket[26]), .Z(n515) );
  N1M2P U302 ( .A(n107), .Z(n307) );
  N1M1P U303 ( .A(n401), .Z(n398) );
  N1M1P U304 ( .A(chosenPacket[28]), .Z(n514) );
  BUFM1P U305 ( .A(N115), .Z(n303) );
  HA1FM1P U306 ( .A(chosenPacket[17]), .B(chosenPacket[16]), .CO(
        \add_x_80_3/carry[2] ), .S(N109) );
  OAI21M2P U307 ( .A(n342), .B(n341), .C(n488), .Z(n349) );
  NR2M1P U308 ( .A(n477), .B(n57), .Z(n473) );
  MUX21LM1P U309 ( .A(Link_Config[0]), .B(Link_Config[2]), .S(N44), .Z(n343)
         );
  MUX21LM1P U310 ( .A(Link_Config[1]), .B(Link_Config[3]), .S(N44), .Z(n342)
         );
  N1M1P U311 ( .A(dataLocation[1]), .Z(n352) );
  ND2BNM1P U312 ( .B(n344), .A(n343), .Z(n348) );
  AOI22M1P U313 ( .A(chosenPacket[21]), .B(n396), .C(n398), .D(N113), .Z(n289)
         );
  AOI22M1P U314 ( .A(Packet_From_Link_W[21]), .B(n320), .C(
        Packet_From_Link_E[21]), .D(n476), .Z(n290) );
  ND3M1P U315 ( .A(n384), .B(n289), .C(n290), .Z(n255) );
  AOI22M1P U316 ( .A(chosenPacket[20]), .B(n396), .C(n398), .D(N112), .Z(n291)
         );
  AOI22M1P U317 ( .A(Packet_From_Link_W[20]), .B(n320), .C(
        Packet_From_Link_E[20]), .D(n476), .Z(n292) );
  ND3M1P U318 ( .A(n385), .B(n291), .C(n292), .Z(n256) );
  AOI22M1P U319 ( .A(chosenPacket[19]), .B(n396), .C(n398), .D(N111), .Z(n293)
         );
  AOI22M1P U320 ( .A(Packet_From_Link_W[19]), .B(n320), .C(
        Packet_From_Link_E[19]), .D(n476), .Z(n294) );
  ND3M1P U321 ( .A(n386), .B(n293), .C(n294), .Z(n257) );
  ND2BNM1P U322 ( .B(Router_Address[7]), .A(chosenPacket[31]), .Z(n367) );
  AOI22M1P U323 ( .A(chosenPacket[18]), .B(n396), .C(n398), .D(N110), .Z(n295)
         );
  AOI22M1P U324 ( .A(Packet_From_Link_W[18]), .B(n320), .C(
        Packet_From_Link_E[18]), .D(n476), .Z(n296) );
  ND3M1P U325 ( .A(n387), .B(n295), .C(n296), .Z(n258) );
  AO211M1P U326 ( .A(n43), .B(Router_Address[5]), .C(n514), .D(
        Router_Address[4]), .Z(n297) );
  AOI22M1P U327 ( .A(n42), .B(Router_Address[6]), .C(n513), .D(n297), .Z(n298)
         );
  ND2BNM1P U328 ( .B(n298), .A(n367), .Z(n299) );
  ND4DNM1P U329 ( .D(TxQueue_Full_E), .A(Link_Config[0]), .B(n369), .C(n299), 
        .Z(n484) );
  NR2BNM1P U330 ( .B(chosenPacket[27]), .A(Router_Address[3]), .Z(n498) );
  AOI22M1P U331 ( .A(Packet_From_Link_E[23]), .B(n306), .C(
        Packet_From_Link_S[23]), .D(n319), .Z(n300) );
  AOI22M1P U332 ( .A(n398), .B(N115), .C(n396), .D(chosenPacket[23]), .Z(n301)
         );
  ND3M1P U333 ( .A(n300), .B(n397), .C(n301), .Z(n262) );
  ND2BNM3P U334 ( .B(n379), .A(n375), .Z(n477) );
  N1M6P U335 ( .A(n311), .Z(n302) );
  N1M3P U336 ( .A(n38), .Z(n311) );
  BUFM8P U337 ( .A(n39), .Z(n333) );
  BUFM6P U338 ( .A(n474), .Z(n318) );
  BUFM4P U339 ( .A(n474), .Z(n319) );
  AND4M1P U340 ( .A(n309), .B(n399), .C(n398), .D(n402), .Z(n40) );
  NR3M2P U341 ( .A(n403), .B(n402), .C(n401), .Z(n39) );
  N1M1P U342 ( .A(chosenPacket[27]), .Z(n44) );
  BUFM2P U343 ( .A(n475), .Z(n320) );
  N1M1P U344 ( .A(n304), .Z(Packet_To_Node[28]) );
  N1M3P U345 ( .A(n400), .Z(n308) );
  NR2FM1P U346 ( .A(n338), .B(n501), .Z(n361) );
  EOFM4P U347 ( .A(\add_x_80_3/carry[7] ), .B(chosenPacket[23]), .Z(N115) );
  HA1M2P U348 ( .A(chosenPacket[20]), .B(\add_x_80_3/carry[4] ), .CO(
        \add_x_80_3/carry[5] ), .S(N112) );
  HA1FM2P U349 ( .A(chosenPacket[21]), .B(\add_x_80_3/carry[5] ), .CO(
        \add_x_80_3/carry[6] ), .S(N113) );
  HA1FM4P U350 ( .A(chosenPacket[22]), .B(\add_x_80_3/carry[6] ), .CO(
        \add_x_80_3/carry[7] ), .S(N114) );
  HA1M2P U351 ( .A(chosenPacket[18]), .B(\add_x_80_3/carry[2] ), .CO(
        \add_x_80_3/carry[3] ), .S(N110) );
  HA1M2P U352 ( .A(chosenPacket[19]), .B(\add_x_80_3/carry[3] ), .CO(
        \add_x_80_3/carry[4] ), .S(N111) );
  NR3M4P U353 ( .A(n482), .B(n334), .C(n484), .Z(n37) );
  N1M6P U354 ( .A(n107), .Z(n329) );
  AOI211M2P U355 ( .A(Router_Address[1]), .B(n45), .C(n494), .D(n498), .Z(n495) );
  N1M8P U356 ( .A(n314), .Z(n316) );
  ND2FM4P U357 ( .A(n488), .B(dataLocation[1]), .Z(n376) );
  AND2M8P U358 ( .A(n339), .B(n6), .Z(n488) );
  N1M6P U359 ( .A(n311), .Z(n312) );
  N1M6P U360 ( .A(n311), .Z(n313) );
  N1M4P U361 ( .A(n314), .Z(n317) );
  N1M4P U362 ( .A(n314), .Z(n315) );
  N1M3P U363 ( .A(n37), .Z(n314) );
  N1M8P U364 ( .A(n308), .Z(n309) );
  N1M8P U365 ( .A(n329), .Z(n327) );
  AOI22M2P U366 ( .A(Router_Address[6]), .B(n42), .C(Router_Address[5]), .D(
        n43), .Z(n508) );
  ND4DNM4P U367 ( .D(TxQueue_Full_N), .A(n365), .B(n507), .C(Link_Config[3]), 
        .Z(n402) );
  N1M4P U368 ( .A(n8), .Z(n490) );
  NR3M3P U369 ( .A(n482), .B(n334), .C(n483), .Z(n38) );
  NR2FM2P U370 ( .A(n477), .B(n6), .Z(n476) );
  AOI22M1P U371 ( .A(RxQueue_Empty_S), .B(n346), .C(RxQueue_Empty_E), .D(n345), 
        .Z(n347) );
  N1M1P U372 ( .A(chosenPacket[25]), .Z(n45) );
  N1M1P U373 ( .A(n486), .Z(n357) );
  ND2FM4P U374 ( .A(n376), .B(n377), .Z(N44) );
  AOI21M4P U375 ( .A(N115), .B(n362), .C(n361), .Z(n400) );
  N1M2P U376 ( .A(n360), .Z(n362) );
  ND4DNFM4P U377 ( .D(n359), .A(N114), .B(N113), .C(N112), .Z(n360) );
  BUFM3P U378 ( .A(n40), .Z(n331) );
  BUFM3P U379 ( .A(n40), .Z(n330) );
  BUFM3P U380 ( .A(n40), .Z(n332) );
  BUFM3P U381 ( .A(n477), .Z(n323) );
  AND2M1P U382 ( .A(n8), .B(Rst_n), .Z(n375) );
  NR2FM1P U383 ( .A(n477), .B(n376), .Z(n478) );
  ND2FM4P U384 ( .A(n340), .B(n352), .Z(n377) );
  NR2M2P U385 ( .A(n510), .B(n493), .Z(n513) );
  N1M4P U386 ( .A(chosenPacket[30]), .Z(n42) );
  ND4DNFM4P U387 ( .D(n399), .A(n309), .B(n490), .C(n402), .Z(n482) );
  NR2FM1P U388 ( .A(n477), .B(n378), .Z(n475) );
  ND4DNFM4P U389 ( .D(n350), .A(n349), .B(n348), .C(n347), .Z(n379) );
  N1M6P U390 ( .A(n329), .Z(n328) );
  OAI22M2P U391 ( .A(Router_Address[2]), .B(n515), .C(Router_Address[1]), .D(
        n45), .Z(n501) );
  N1M2P U392 ( .A(chosenPacket[24]), .Z(n492) );
  N1M2P U393 ( .A(chosenPacket[29]), .Z(n43) );
  BUFM2P U394 ( .A(n475), .Z(n322) );
  BUFM2P U395 ( .A(n475), .Z(n321) );
  ND2M2P U396 ( .A(n340), .B(dataLocation[1]), .Z(n57) );
  AND2M2P U397 ( .A(n361), .B(n490), .Z(n489) );
  ND2M1P U398 ( .A(n490), .B(Rst_n), .Z(n401) );
  N1M1P U399 ( .A(dataLocation[0]), .Z(n339) );
  N1M1P U400 ( .A(Rst_n), .Z(n334) );
  AOI21M1P U401 ( .A(n506), .B(n507), .C(n358), .Z(n399) );
  ND2M1P U402 ( .A(Router_Address[3]), .B(n44), .Z(n507) );
  N1M1P U403 ( .A(chosenPacket[31]), .Z(n491) );
  OAI22M1P U404 ( .A(n357), .B(n57), .C(n490), .D(n356), .Z(n245) );
  N1M1P U405 ( .A(Node_Read), .Z(n356) );
  OAI22M1P U406 ( .A(n357), .B(n378), .C(n490), .D(n353), .Z(n248) );
  N1M1P U407 ( .A(RxQueue_Read_W), .Z(n353) );
  OAI22M1P U408 ( .A(n357), .B(n376), .C(n490), .D(n355), .Z(n246) );
  N1M1P U409 ( .A(RxQueue_Read_N), .Z(n355) );
  OAI22M1P U410 ( .A(n357), .B(n6), .C(n351), .D(n490), .Z(n249) );
  N1M1P U411 ( .A(RxQueue_Read_E), .Z(n351) );
  OAI22M1P U412 ( .A(n357), .B(n377), .C(n490), .D(n354), .Z(n247) );
  N1M1P U413 ( .A(RxQueue_Read_S), .Z(n354) );
  AOI21M1P U414 ( .A(n372), .B(n371), .C(n8), .Z(n252) );
  N1M1P U415 ( .A(TxQueue_Write_S), .Z(n371) );
  ND3M1P U416 ( .A(n309), .B(n399), .C(n402), .Z(n372) );
  NR2M1P U417 ( .A(n374), .B(n8), .Z(n253) );
  AOI21M1P U418 ( .A(n309), .B(n373), .C(TxQueue_Write_N), .Z(n374) );
  N1M1P U419 ( .A(n402), .Z(n373) );
  AOI22M1P U420 ( .A(n324), .B(Packet_From_Link_N[21]), .C(n474), .D(
        Packet_From_Link_S[21]), .Z(n384) );
  AOI22M1P U421 ( .A(n324), .B(Packet_From_Link_N[18]), .C(n319), .D(
        Packet_From_Link_S[18]), .Z(n387) );
  AOI22M1P U422 ( .A(n324), .B(Packet_From_Link_N[19]), .C(n319), .D(
        Packet_From_Link_S[19]), .Z(n386) );
  AOI22M1P U423 ( .A(n324), .B(Packet_From_Link_N[20]), .C(n319), .D(
        Packet_From_Link_S[20]), .Z(n385) );
  ND4M1P U424 ( .A(n395), .B(n394), .C(n393), .D(n392), .Z(n260) );
  MUX21LM1P U425 ( .A(n398), .B(n396), .S(chosenPacket[16]), .Z(n392) );
  ND2M1P U426 ( .A(n476), .B(Packet_From_Link_E[16]), .Z(n393) );
  ND2M1P U427 ( .A(n320), .B(Packet_From_Link_W[16]), .Z(n394) );
  AOI22M1P U428 ( .A(n324), .B(Packet_From_Link_N[16]), .C(n319), .D(
        Packet_From_Link_S[16]), .Z(n395) );
  OAI22M1P U429 ( .A(n482), .B(n484), .C(n8), .D(n366), .Z(n250) );
  N1M1P U430 ( .A(TxQueue_Write_E), .Z(n366) );
  OAI22M1P U431 ( .A(n482), .B(n483), .C(n8), .D(n370), .Z(n251) );
  N1M1P U432 ( .A(TxQueue_Write_W), .Z(n370) );
  ND4M1P U433 ( .A(n383), .B(n382), .C(n381), .D(n380), .Z(n254) );
  ND2M1P U434 ( .A(n476), .B(Packet_From_Link_E[22]), .Z(n381) );
  ND2M1P U435 ( .A(n320), .B(Packet_From_Link_W[22]), .Z(n382) );
  AOI22M1P U436 ( .A(n324), .B(Packet_From_Link_N[22]), .C(n474), .D(
        Packet_From_Link_S[22]), .Z(n383) );
  ND2M1P U437 ( .A(n476), .B(Packet_From_Link_E[17]), .Z(n389) );
  ND2M1P U438 ( .A(n320), .B(Packet_From_Link_W[17]), .Z(n390) );
  AOI22M1P U439 ( .A(n324), .B(Packet_From_Link_N[17]), .C(n319), .D(
        Packet_From_Link_S[17]), .Z(n391) );
  AOI211M1P U440 ( .A(n489), .B(To_Node_Full), .C(n487), .D(n486), .Z(n7) );
  NR2M1P U441 ( .A(n379), .B(n490), .Z(n486) );
  AND3M1P U442 ( .A(n485), .B(n484), .C(n483), .Z(n487) );
  N1M1P U443 ( .A(n309), .Z(n403) );
  ND3M1P U444 ( .A(n457), .B(n456), .C(n455), .Z(n269) );
  AOI22M1P U445 ( .A(Packet_From_Link_N[25]), .B(n326), .C(chosenPacket[25]), 
        .D(n323), .Z(n455) );
  AOI22M1P U446 ( .A(n306), .B(Packet_From_Link_E[25]), .C(n321), .D(
        Packet_From_Link_W[25]), .Z(n456) );
  AOI22M1P U447 ( .A(n318), .B(Packet_From_Link_S[25]), .C(n305), .D(
        Packet_From_Node_25), .Z(n457) );
  ND3M1P U448 ( .A(n469), .B(n468), .C(n467), .Z(n265) );
  AOI22M1P U449 ( .A(Packet_From_Link_N[29]), .B(n326), .C(chosenPacket[29]), 
        .D(n323), .Z(n467) );
  AOI22M1P U450 ( .A(n306), .B(Packet_From_Link_E[29]), .C(n321), .D(
        Packet_From_Link_W[29]), .Z(n468) );
  AOI22M1P U451 ( .A(n318), .B(Packet_From_Link_S[29]), .C(n305), .D(
        Packet_From_Node_29), .Z(n469) );
  ND3M1P U452 ( .A(n454), .B(n453), .C(n452), .Z(n270) );
  AOI22M1P U453 ( .A(Packet_From_Link_N[24]), .B(n326), .C(chosenPacket[24]), 
        .D(n323), .Z(n452) );
  AOI22M1P U454 ( .A(n306), .B(Packet_From_Link_E[24]), .C(n321), .D(
        Packet_From_Link_W[24]), .Z(n453) );
  AOI22M1P U455 ( .A(n318), .B(Packet_From_Link_S[24]), .C(n305), .D(
        Packet_From_Node_24), .Z(n454) );
  AO21CNM1P U456 ( .A(n379), .B(n8), .C(Rst_n), .Z(n396) );
  AOI22M1P U457 ( .A(n324), .B(Packet_From_Link_N[23]), .C(n320), .D(
        Packet_From_Link_W[23]), .Z(n397) );
  ND3M1P U458 ( .A(n415), .B(n414), .C(n413), .Z(n283) );
  AOI22M1P U459 ( .A(Packet_From_Link_N[3]), .B(n325), .C(chosenPacket[3]), 
        .D(n323), .Z(n413) );
  AOI22M1P U460 ( .A(n306), .B(Packet_From_Link_E[3]), .C(n320), .D(
        Packet_From_Link_W[3]), .Z(n414) );
  AOI22M1P U461 ( .A(n319), .B(Packet_From_Link_S[3]), .C(n305), .D(
        Packet_From_Node[3]), .Z(n415) );
  ND3M1P U462 ( .A(n412), .B(n411), .C(n410), .Z(n284) );
  AOI22M1P U463 ( .A(Packet_From_Link_N[2]), .B(n325), .C(chosenPacket[2]), 
        .D(n323), .Z(n410) );
  AOI22M1P U464 ( .A(n306), .B(Packet_From_Link_E[2]), .C(n320), .D(
        Packet_From_Link_W[2]), .Z(n411) );
  AOI22M1P U465 ( .A(n319), .B(Packet_From_Link_S[2]), .C(n305), .D(
        Packet_From_Node[2]), .Z(n412) );
  ND3M1P U466 ( .A(n409), .B(n408), .C(n407), .Z(n285) );
  AOI22M1P U467 ( .A(Packet_From_Link_N[1]), .B(n324), .C(chosenPacket[1]), 
        .D(n323), .Z(n407) );
  AOI22M1P U468 ( .A(n306), .B(Packet_From_Link_E[1]), .C(n320), .D(
        Packet_From_Link_W[1]), .Z(n408) );
  AOI22M1P U469 ( .A(n319), .B(Packet_From_Link_S[1]), .C(n305), .D(
        Packet_From_Node[1]), .Z(n409) );
  ND3M1P U470 ( .A(n406), .B(n405), .C(n404), .Z(n286) );
  AOI22M1P U471 ( .A(Packet_From_Link_N[0]), .B(n324), .C(chosenPacket[0]), 
        .D(n323), .Z(n404) );
  AOI22M1P U472 ( .A(n306), .B(Packet_From_Link_E[0]), .C(n320), .D(
        Packet_From_Link_W[0]), .Z(n405) );
  AOI22M1P U473 ( .A(n319), .B(Packet_From_Link_S[0]), .C(n305), .D(
        Packet_From_Node[0]), .Z(n406) );
  ND3M1P U474 ( .A(n430), .B(n429), .C(n428), .Z(n278) );
  AOI22M1P U475 ( .A(Packet_From_Link_N[8]), .B(n325), .C(chosenPacket[8]), 
        .D(n323), .Z(n428) );
  AOI22M1P U476 ( .A(n306), .B(Packet_From_Link_E[8]), .C(n322), .D(
        Packet_From_Link_W[8]), .Z(n429) );
  AOI22M1P U477 ( .A(n318), .B(Packet_From_Link_S[8]), .C(n305), .D(
        Packet_From_Node[8]), .Z(n430) );
  ND3M1P U478 ( .A(n472), .B(n471), .C(n470), .Z(n264) );
  AOI22M1P U479 ( .A(Packet_From_Link_N[30]), .B(n478), .C(chosenPacket[30]), 
        .D(n323), .Z(n470) );
  AOI22M1P U480 ( .A(n306), .B(Packet_From_Link_E[30]), .C(n321), .D(
        Packet_From_Link_W[30]), .Z(n471) );
  AOI22M1P U481 ( .A(n318), .B(Packet_From_Link_S[30]), .C(n305), .D(
        Packet_From_Node_30), .Z(n472) );
  ND3M1P U482 ( .A(n451), .B(n450), .C(n449), .Z(n271) );
  AOI22M1P U483 ( .A(Packet_From_Link_N[15]), .B(n326), .C(chosenPacket[15]), 
        .D(n323), .Z(n449) );
  AOI22M1P U484 ( .A(n306), .B(Packet_From_Link_E[15]), .C(n321), .D(
        Packet_From_Link_W[15]), .Z(n450) );
  AOI22M1P U485 ( .A(n318), .B(Packet_From_Link_S[15]), .C(n305), .D(
        Packet_From_Node[15]), .Z(n451) );
  ND3M1P U486 ( .A(n463), .B(n462), .C(n461), .Z(n267) );
  AOI22M1P U487 ( .A(Packet_From_Link_N[27]), .B(n326), .C(chosenPacket[27]), 
        .D(n323), .Z(n461) );
  AOI22M1P U488 ( .A(n306), .B(Packet_From_Link_E[27]), .C(n321), .D(
        Packet_From_Link_W[27]), .Z(n462) );
  AOI22M1P U489 ( .A(n318), .B(Packet_From_Link_S[27]), .C(n305), .D(
        Packet_From_Node_27), .Z(n463) );
  ND3M1P U490 ( .A(n427), .B(n426), .C(n425), .Z(n279) );
  AOI22M1P U491 ( .A(Packet_From_Link_N[7]), .B(n325), .C(chosenPacket[7]), 
        .D(n323), .Z(n425) );
  AOI22M1P U492 ( .A(n306), .B(Packet_From_Link_E[7]), .C(n322), .D(
        Packet_From_Link_W[7]), .Z(n426) );
  AOI22M1P U493 ( .A(n318), .B(Packet_From_Link_S[7]), .C(n305), .D(
        Packet_From_Node[7]), .Z(n427) );
  ND3M1P U494 ( .A(n448), .B(n447), .C(n446), .Z(n272) );
  AOI22M1P U495 ( .A(Packet_From_Link_N[14]), .B(n326), .C(chosenPacket[14]), 
        .D(n323), .Z(n446) );
  AOI22M1P U496 ( .A(n306), .B(Packet_From_Link_E[14]), .C(n321), .D(
        Packet_From_Link_W[14]), .Z(n447) );
  AOI22M1P U497 ( .A(n318), .B(Packet_From_Link_S[14]), .C(n305), .D(
        Packet_From_Node[14]), .Z(n448) );
  ND3M1P U498 ( .A(n418), .B(n417), .C(n416), .Z(n282) );
  AOI22M1P U499 ( .A(Packet_From_Link_N[4]), .B(n325), .C(chosenPacket[4]), 
        .D(n323), .Z(n416) );
  AOI22M1P U500 ( .A(n306), .B(Packet_From_Link_E[4]), .C(n322), .D(
        Packet_From_Link_W[4]), .Z(n417) );
  AOI22M1P U501 ( .A(n319), .B(Packet_From_Link_S[4]), .C(n305), .D(
        Packet_From_Node[4]), .Z(n418) );
  ND3M1P U502 ( .A(n445), .B(n444), .C(n443), .Z(n273) );
  AOI22M1P U503 ( .A(Packet_From_Link_N[13]), .B(n326), .C(chosenPacket[13]), 
        .D(n323), .Z(n443) );
  AOI22M1P U504 ( .A(n306), .B(Packet_From_Link_E[13]), .C(n322), .D(
        Packet_From_Link_W[13]), .Z(n444) );
  AOI22M1P U505 ( .A(n318), .B(Packet_From_Link_S[13]), .C(n305), .D(
        Packet_From_Node[13]), .Z(n445) );
  ND3M1P U506 ( .A(n433), .B(n432), .C(n431), .Z(n277) );
  AOI22M1P U507 ( .A(Packet_From_Link_N[9]), .B(n325), .C(chosenPacket[9]), 
        .D(n323), .Z(n431) );
  AOI22M1P U508 ( .A(n306), .B(Packet_From_Link_E[9]), .C(n322), .D(
        Packet_From_Link_W[9]), .Z(n432) );
  AOI22M1P U509 ( .A(n319), .B(Packet_From_Link_S[9]), .C(n305), .D(
        Packet_From_Node[9]), .Z(n433) );
  ND3M1P U510 ( .A(n421), .B(n420), .C(n419), .Z(n281) );
  AOI22M1P U511 ( .A(Packet_From_Link_N[5]), .B(n325), .C(chosenPacket[5]), 
        .D(n323), .Z(n419) );
  AOI22M1P U512 ( .A(n306), .B(Packet_From_Link_E[5]), .C(n322), .D(
        Packet_From_Link_W[5]), .Z(n420) );
  AOI22M1P U513 ( .A(n318), .B(Packet_From_Link_S[5]), .C(n305), .D(
        Packet_From_Node[5]), .Z(n421) );
  ND3M1P U514 ( .A(n442), .B(n441), .C(n440), .Z(n274) );
  AOI22M1P U515 ( .A(Packet_From_Link_N[12]), .B(n326), .C(chosenPacket[12]), 
        .D(n323), .Z(n440) );
  AOI22M1P U516 ( .A(n306), .B(Packet_From_Link_E[12]), .C(n322), .D(
        Packet_From_Link_W[12]), .Z(n441) );
  AOI22M1P U517 ( .A(n319), .B(Packet_From_Link_S[12]), .C(n305), .D(
        Packet_From_Node[12]), .Z(n442) );
  ND3M1P U518 ( .A(n424), .B(n423), .C(n422), .Z(n280) );
  AOI22M1P U519 ( .A(Packet_From_Link_N[6]), .B(n325), .C(chosenPacket[6]), 
        .D(n323), .Z(n422) );
  AOI22M1P U520 ( .A(n306), .B(Packet_From_Link_E[6]), .C(n322), .D(
        Packet_From_Link_W[6]), .Z(n423) );
  AOI22M1P U521 ( .A(n318), .B(Packet_From_Link_S[6]), .C(n305), .D(
        Packet_From_Node[6]), .Z(n424) );
  ND3M1P U522 ( .A(n439), .B(n438), .C(n437), .Z(n275) );
  AOI22M1P U523 ( .A(Packet_From_Link_N[11]), .B(n325), .C(chosenPacket[11]), 
        .D(n323), .Z(n437) );
  AOI22M1P U524 ( .A(n306), .B(Packet_From_Link_E[11]), .C(n322), .D(
        Packet_From_Link_W[11]), .Z(n438) );
  AOI22M1P U525 ( .A(n319), .B(Packet_From_Link_S[11]), .C(n305), .D(
        Packet_From_Node[11]), .Z(n439) );
  ND3M1P U526 ( .A(n436), .B(n435), .C(n434), .Z(n276) );
  AOI22M1P U527 ( .A(Packet_From_Link_N[10]), .B(n325), .C(chosenPacket[10]), 
        .D(n323), .Z(n434) );
  AOI22M1P U528 ( .A(n306), .B(Packet_From_Link_E[10]), .C(n322), .D(
        Packet_From_Link_W[10]), .Z(n435) );
  AOI22M1P U529 ( .A(n318), .B(Packet_From_Link_S[10]), .C(n305), .D(
        Packet_From_Node[10]), .Z(n436) );
  ND3M1P U530 ( .A(n481), .B(n480), .C(n479), .Z(n263) );
  AOI22M1P U531 ( .A(Packet_From_Link_N[31]), .B(n478), .C(chosenPacket[31]), 
        .D(n323), .Z(n479) );
  AOI22M1P U532 ( .A(n306), .B(Packet_From_Link_E[31]), .C(n321), .D(
        Packet_From_Link_W[31]), .Z(n480) );
  AOI22M1P U533 ( .A(n318), .B(Packet_From_Link_S[31]), .C(n305), .D(
        Packet_From_Node_31), .Z(n481) );
  ND3M1P U534 ( .A(n460), .B(n459), .C(n458), .Z(n268) );
  AOI22M1P U535 ( .A(Packet_From_Link_N[26]), .B(n326), .C(chosenPacket[26]), 
        .D(n323), .Z(n458) );
  AOI22M1P U536 ( .A(n306), .B(Packet_From_Link_E[26]), .C(n321), .D(
        Packet_From_Link_W[26]), .Z(n459) );
  AOI22M1P U537 ( .A(n318), .B(Packet_From_Link_S[26]), .C(n305), .D(
        Packet_From_Node_26), .Z(n460) );
  ND3M1P U538 ( .A(n466), .B(n465), .C(n464), .Z(n266) );
  AOI22M1P U539 ( .A(Packet_From_Link_N[28]), .B(n326), .C(chosenPacket[28]), 
        .D(n323), .Z(n464) );
  AOI22M1P U540 ( .A(n306), .B(Packet_From_Link_E[28]), .C(n321), .D(
        Packet_From_Link_W[28]), .Z(n465) );
  ND2M1P U541 ( .A(n488), .B(n352), .Z(n378) );
  AOI22M1P U542 ( .A(n318), .B(Packet_From_Link_S[28]), .C(n305), .D(
        Packet_From_Node_28), .Z(n466) );
  N1M1P U543 ( .A(n6), .Z(n345) );
  N1M1P U544 ( .A(n377), .Z(n346) );
  ND2BNM1P U545 ( .B(n488), .A(n57), .Z(n344) );
  MUX21HM1P U546 ( .A(RxQueue_Empty_W), .B(RxQueue_Empty_N), .S(
        dataLocation[1]), .Z(n341) );
  NR2BNM1P U547 ( .B(Node_Queue_Empty), .A(n57), .Z(n350) );
  ND2BNM1P U548 ( .B(chosenPacket[31]), .A(Router_Address[7]), .Z(n369) );
  OAI21M1P U549 ( .A(n364), .B(n505), .C(n363), .Z(n365) );
  N1M1P U550 ( .A(n498), .Z(n363) );
  NR2M1P U551 ( .A(n501), .B(n499), .Z(n364) );
  ND4M1P U552 ( .A(N111), .B(N110), .C(N109), .D(n310), .Z(n359) );
  ND2BNM1P U553 ( .B(TxQueue_Full_S), .A(Link_Config[2]), .Z(n358) );
  NR2BNM4P U554 ( .B(n489), .A(To_Node_Full), .Z(n107) );
  ENFM1P U555 ( .A(Router_Address[7]), .B(chosenPacket[31]), .Z(n335) );
  N1M1P U556 ( .A(Router_Address[0]), .Z(n336) );
  ND4M1P U557 ( .A(n513), .B(n508), .C(n495), .D(n500), .Z(n496) );
  NR2M1P U558 ( .A(Router_Address[0]), .B(n492), .Z(n494) );
  MUX21HM1P U559 ( .A(Packet_To_Node[18]), .B(N110), .S(n328), .Z(n27) );
  MUX21HM1P U560 ( .A(Packet_To_Node[19]), .B(N111), .S(n327), .Z(n28) );
  MUX21HM1P U561 ( .A(Packet_To_Node[20]), .B(N112), .S(n328), .Z(n29) );
  MUX21HM1P U562 ( .A(Packet_To_Node[21]), .B(N113), .S(n328), .Z(n30) );
  MUX21HM1P U563 ( .A(Packet_To_Node[17]), .B(N109), .S(n328), .Z(n26) );
  N1M1P U564 ( .A(chosenPacket[16]), .Z(n310) );
  OAI211M1P U565 ( .A(Router_Address[4]), .B(n514), .C(n507), .D(n509), .Z(
        n497) );
  ND4M1P U566 ( .A(n391), .B(n390), .C(n389), .D(n388), .Z(n259) );
  MUX21HM1P U567 ( .A(Packet_To_Node[23]), .B(N115), .S(n328), .Z(n32) );
  AOI22M1P U568 ( .A(chosenPacket[22]), .B(n396), .C(N114), .D(n398), .Z(n380)
         );
  AOI22M1P U569 ( .A(chosenPacket[17]), .B(n396), .C(N109), .D(n398), .Z(n388)
         );
  N1M1P U570 ( .A(n482), .Z(n485) );
  OAI21M1P U571 ( .A(chosenPacket[24]), .B(n336), .C(n335), .Z(n337) );
  OR3M1P U572 ( .A(n496), .B(n497), .C(n337), .Z(n338) );
  MUX21HM1P U573 ( .A(Packet_To_Node[22]), .B(N114), .S(n328), .Z(n31) );
  ND3CNM1P U574 ( .C(TxQueue_Full_W), .A(n367), .B(Link_Config[1]), .Z(n368)
         );
  AO21M1P U575 ( .A(n512), .B(n369), .C(n368), .Z(n483) );
  ND2M1P U576 ( .A(Router_Address[4]), .B(n514), .Z(n509) );
  NR2M1P U577 ( .A(Router_Address[5]), .B(n43), .Z(n510) );
  NR2M1P U578 ( .A(Router_Address[6]), .B(n42), .Z(n493) );
  ND2M1P U579 ( .A(Router_Address[2]), .B(n515), .Z(n500) );
  AO21CNM1P U580 ( .A(To_Node_Write), .B(n490), .C(n307), .Z(n261) );
  AOI211M1P U581 ( .A(Router_Address[1]), .B(n45), .C(Router_Address[0]), .D(
        n492), .Z(n499) );
  N1M1P U582 ( .A(n500), .Z(n505) );
  ND2M1P U583 ( .A(Router_Address[1]), .B(n45), .Z(n503) );
  ND2M1P U584 ( .A(Router_Address[0]), .B(n492), .Z(n502) );
  AOI21M1P U585 ( .A(n503), .B(n502), .C(n501), .Z(n504) );
  OAI22M1P U586 ( .A(Router_Address[3]), .B(n44), .C(n505), .D(n504), .Z(n506)
         );
  OAI21M1P U587 ( .A(n510), .B(n509), .C(n508), .Z(n511) );
  OAI21M1P U588 ( .A(Router_Address[6]), .B(n42), .C(n511), .Z(n512) );
  AOI22DNM1P U589 ( .A(n327), .B(n515), .D(Packet_To_Node[26]), .C(n329), .Z(
        n34) );
  AOI22DNM1P U590 ( .A(n327), .B(n492), .D(Packet_To_Node[24]), .C(n329), .Z(
        n33) );
  AOI22DNM1P U591 ( .A(n327), .B(chosenPacket[16]), .D(Packet_To_Node[16]), 
        .C(n329), .Z(n25) );
  OAI22M1P U592 ( .A(n307), .B(chosenPacket[15]), .C(Packet_To_Node[15]), .D(
        n328), .Z(n516) );
  N1M1P U593 ( .A(n516), .Z(n24) );
  OAI22M1P U594 ( .A(n307), .B(chosenPacket[14]), .C(Packet_To_Node[14]), .D(
        n327), .Z(n517) );
  N1M1P U595 ( .A(n517), .Z(n23) );
  OAI22M1P U596 ( .A(n307), .B(chosenPacket[13]), .C(Packet_To_Node[13]), .D(
        n328), .Z(n518) );
  N1M1P U597 ( .A(n518), .Z(n22) );
  OAI22M1P U598 ( .A(n307), .B(chosenPacket[12]), .C(Packet_To_Node[12]), .D(
        n327), .Z(n519) );
  N1M1P U599 ( .A(n519), .Z(n21) );
  OAI22M1P U600 ( .A(n307), .B(chosenPacket[11]), .C(Packet_To_Node[11]), .D(
        n327), .Z(n520) );
  N1M1P U601 ( .A(n520), .Z(n20) );
  OAI22M1P U602 ( .A(n307), .B(chosenPacket[10]), .C(Packet_To_Node[10]), .D(
        n327), .Z(n521) );
  N1M1P U603 ( .A(n521), .Z(n19) );
  OAI22M1P U604 ( .A(n307), .B(chosenPacket[9]), .C(Packet_To_Node[9]), .D(
        n327), .Z(n522) );
  N1M1P U605 ( .A(n522), .Z(n18) );
  OAI22M1P U606 ( .A(n307), .B(chosenPacket[8]), .C(Packet_To_Node[8]), .D(
        n327), .Z(n523) );
  N1M1P U607 ( .A(n523), .Z(n17) );
  OAI22M1P U608 ( .A(n307), .B(chosenPacket[7]), .C(Packet_To_Node[7]), .D(
        n327), .Z(n524) );
  N1M1P U609 ( .A(n524), .Z(n16) );
  OAI22M1P U610 ( .A(n307), .B(chosenPacket[6]), .C(Packet_To_Node[6]), .D(
        n328), .Z(n525) );
  N1M1P U611 ( .A(n525), .Z(n15) );
  OAI22M1P U612 ( .A(n307), .B(chosenPacket[5]), .C(Packet_To_Node[5]), .D(
        n328), .Z(n526) );
  N1M1P U613 ( .A(n526), .Z(n14) );
  OAI22M1P U614 ( .A(n307), .B(chosenPacket[4]), .C(Packet_To_Node[4]), .D(
        n328), .Z(n527) );
  N1M1P U615 ( .A(n527), .Z(n13) );
  OAI22M1P U616 ( .A(n307), .B(chosenPacket[3]), .C(Packet_To_Node[3]), .D(
        n328), .Z(n528) );
  N1M1P U617 ( .A(n528), .Z(n12) );
  OAI22M1P U618 ( .A(n307), .B(chosenPacket[2]), .C(Packet_To_Node[2]), .D(
        n328), .Z(n529) );
  N1M1P U619 ( .A(n529), .Z(n11) );
  OAI22M1P U620 ( .A(n307), .B(chosenPacket[1]), .C(Packet_To_Node[1]), .D(
        n328), .Z(n530) );
  N1M1P U621 ( .A(n530), .Z(n10) );
  OAI22M1P U622 ( .A(n307), .B(chosenPacket[0]), .C(Packet_To_Node[0]), .D(
        n328), .Z(n531) );
  N1M1P U623 ( .A(n531), .Z(n9) );
  N1M1P U624 ( .A(n5), .Z(Packet_To_Node[31]) );
  N1M1P U625 ( .A(n4), .Z(Packet_To_Node[30]) );
  N1M1P U626 ( .A(n3), .Z(Packet_To_Node[29]) );
  N1M1P U627 ( .A(n2), .Z(Packet_To_Node[27]) );
  N1M1P U628 ( .A(n1), .Z(Packet_To_Node[25]) );
endmodule

