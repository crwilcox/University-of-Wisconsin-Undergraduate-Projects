library verilog;
use verilog.vl_types.all;
entity decoder_2_to_4_139_tb is
end decoder_2_to_4_139_tb;
