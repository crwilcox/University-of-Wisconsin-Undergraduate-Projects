library verilog;
use verilog.vl_types.all;
entity partial_counter_tb is
end partial_counter_tb;
