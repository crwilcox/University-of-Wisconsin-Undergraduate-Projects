library verilog;
use verilog.vl_types.all;
entity prime_detector_structural_tb is
end prime_detector_structural_tb;
