
module Packet_Queue_0 ( Clk_r, Rst_n, Packet_In, Read_Ack, Write_Ack, 
        Packet_Out, Empty, Full );
  input [31:0] Packet_In;
  output [31:0] Packet_Out;
  input Clk_r, Rst_n, Read_Ack, Write_Ack;
  output Empty, Full;
  wire   \Queue[4][31] , \Queue[4][30] , \Queue[4][29] , \Queue[4][28] ,
         \Queue[4][27] , \Queue[4][26] , \Queue[4][25] , \Queue[4][24] ,
         \Queue[4][23] , \Queue[4][22] , \Queue[4][21] , \Queue[4][20] ,
         \Queue[4][19] , \Queue[4][18] , \Queue[4][17] , \Queue[4][16] ,
         \Queue[4][15] , \Queue[4][14] , \Queue[4][13] , \Queue[4][12] ,
         \Queue[4][11] , \Queue[4][10] , \Queue[4][9] , \Queue[4][8] ,
         \Queue[4][7] , \Queue[4][6] , \Queue[4][5] , \Queue[4][4] ,
         \Queue[4][3] , \Queue[4][2] , \Queue[4][1] , \Queue[4][0] ,
         \Queue[3][31] , \Queue[3][30] , \Queue[3][29] , \Queue[3][28] ,
         \Queue[3][27] , \Queue[3][26] , \Queue[3][25] , \Queue[3][24] ,
         \Queue[3][23] , \Queue[3][22] , \Queue[3][21] , \Queue[3][20] ,
         \Queue[3][19] , \Queue[3][18] , \Queue[3][17] , \Queue[3][16] ,
         \Queue[3][15] , \Queue[3][14] , \Queue[3][13] , \Queue[3][12] ,
         \Queue[3][11] , \Queue[3][10] , \Queue[3][9] , \Queue[3][8] ,
         \Queue[3][7] , \Queue[3][6] , \Queue[3][5] , \Queue[3][4] ,
         \Queue[3][3] , \Queue[3][2] , \Queue[3][1] , \Queue[3][0] ,
         \Queue[2][31] , \Queue[2][30] , \Queue[2][29] , \Queue[2][28] ,
         \Queue[2][27] , \Queue[2][26] , \Queue[2][25] , \Queue[2][24] ,
         \Queue[2][23] , \Queue[2][22] , \Queue[2][21] , \Queue[2][20] ,
         \Queue[2][19] , \Queue[2][18] , \Queue[2][17] , \Queue[2][16] ,
         \Queue[2][15] , \Queue[2][14] , \Queue[2][13] , \Queue[2][12] ,
         \Queue[2][11] , \Queue[2][10] , \Queue[2][9] , \Queue[2][8] ,
         \Queue[2][7] , \Queue[2][6] , \Queue[2][5] , \Queue[2][4] ,
         \Queue[2][3] , \Queue[2][2] , \Queue[2][1] , \Queue[2][0] ,
         \Queue[1][31] , \Queue[1][30] , \Queue[1][29] , \Queue[1][28] ,
         \Queue[1][27] , \Queue[1][26] , \Queue[1][25] , \Queue[1][24] ,
         \Queue[1][23] , \Queue[1][22] , \Queue[1][21] , \Queue[1][20] ,
         \Queue[1][19] , \Queue[1][18] , \Queue[1][17] , \Queue[1][16] ,
         \Queue[1][15] , \Queue[1][14] , \Queue[1][13] , \Queue[1][12] ,
         \Queue[1][11] , \Queue[1][10] , \Queue[1][9] , \Queue[1][8] ,
         \Queue[1][7] , \Queue[1][6] , \Queue[1][5] , \Queue[1][4] ,
         \Queue[1][3] , \Queue[1][2] , \Queue[1][1] , \Queue[1][0] , n1, n2,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n373, n374, n375, n376;
  wire   [2:0] Count;

  FDN2QM1P \Count_reg[0]  ( .D(n372), .CPN(Clk_r), .CD(Rst_n), .Q(Count[0]) );
  FDN2QM1P \Count_reg[1]  ( .D(n371), .CPN(Clk_r), .CD(Rst_n), .Q(Count[1]) );
  FDN2QM1P \Count_reg[2]  ( .D(n370), .CPN(Clk_r), .CD(Rst_n), .Q(Count[2]) );
  FDN1QM1P \Queue_reg[4][30]  ( .D(n338), .CPN(Clk_r), .Q(\Queue[4][30] ) );
  FDN1QM1P \Queue_reg[3][30]  ( .D(n210), .CPN(Clk_r), .Q(\Queue[3][30] ) );
  FDN1QM1P \Queue_reg[2][30]  ( .D(n242), .CPN(Clk_r), .Q(\Queue[2][30] ) );
  FDN1QM1P \Queue_reg[4][29]  ( .D(n339), .CPN(Clk_r), .Q(\Queue[4][29] ) );
  FDN1QM1P \Queue_reg[3][29]  ( .D(n211), .CPN(Clk_r), .Q(\Queue[3][29] ) );
  FDN1QM1P \Queue_reg[2][29]  ( .D(n243), .CPN(Clk_r), .Q(\Queue[2][29] ) );
  FDN1QM1P \Queue_reg[4][28]  ( .D(n340), .CPN(Clk_r), .Q(\Queue[4][28] ) );
  FDN1QM1P \Queue_reg[3][28]  ( .D(n212), .CPN(Clk_r), .Q(\Queue[3][28] ) );
  FDN1QM1P \Queue_reg[2][28]  ( .D(n244), .CPN(Clk_r), .Q(\Queue[2][28] ) );
  FDN1QM1P \Queue_reg[4][27]  ( .D(n341), .CPN(Clk_r), .Q(\Queue[4][27] ) );
  FDN1QM1P \Queue_reg[3][27]  ( .D(n213), .CPN(Clk_r), .Q(\Queue[3][27] ) );
  FDN1QM1P \Queue_reg[2][27]  ( .D(n245), .CPN(Clk_r), .Q(\Queue[2][27] ) );
  FDN1QM1P \Queue_reg[4][26]  ( .D(n342), .CPN(Clk_r), .Q(\Queue[4][26] ) );
  FDN1QM1P \Queue_reg[3][26]  ( .D(n214), .CPN(Clk_r), .Q(\Queue[3][26] ) );
  FDN1QM1P \Queue_reg[2][26]  ( .D(n246), .CPN(Clk_r), .Q(\Queue[2][26] ) );
  FDN1QM1P \Queue_reg[4][25]  ( .D(n343), .CPN(Clk_r), .Q(\Queue[4][25] ) );
  FDN1QM1P \Queue_reg[3][25]  ( .D(n215), .CPN(Clk_r), .Q(\Queue[3][25] ) );
  FDN1QM1P \Queue_reg[2][25]  ( .D(n247), .CPN(Clk_r), .Q(\Queue[2][25] ) );
  FDN1QM1P \Queue_reg[4][24]  ( .D(n344), .CPN(Clk_r), .Q(\Queue[4][24] ) );
  FDN1QM1P \Queue_reg[3][24]  ( .D(n216), .CPN(Clk_r), .Q(\Queue[3][24] ) );
  FDN1QM1P \Queue_reg[2][24]  ( .D(n248), .CPN(Clk_r), .Q(\Queue[2][24] ) );
  FDN1QM1P \Queue_reg[4][23]  ( .D(n345), .CPN(Clk_r), .Q(\Queue[4][23] ) );
  FDN1QM1P \Queue_reg[3][23]  ( .D(n217), .CPN(Clk_r), .Q(\Queue[3][23] ) );
  FDN1QM1P \Queue_reg[2][23]  ( .D(n249), .CPN(Clk_r), .Q(\Queue[2][23] ) );
  FDN1QM1P \Queue_reg[4][22]  ( .D(n346), .CPN(Clk_r), .Q(\Queue[4][22] ) );
  FDN1QM1P \Queue_reg[3][22]  ( .D(n218), .CPN(Clk_r), .Q(\Queue[3][22] ) );
  FDN1QM1P \Queue_reg[2][22]  ( .D(n250), .CPN(Clk_r), .Q(\Queue[2][22] ) );
  FDN1QM1P \Queue_reg[4][21]  ( .D(n347), .CPN(Clk_r), .Q(\Queue[4][21] ) );
  FDN1QM1P \Queue_reg[3][21]  ( .D(n219), .CPN(Clk_r), .Q(\Queue[3][21] ) );
  FDN1QM1P \Queue_reg[2][21]  ( .D(n251), .CPN(Clk_r), .Q(\Queue[2][21] ) );
  FDN1QM1P \Queue_reg[4][20]  ( .D(n348), .CPN(Clk_r), .Q(\Queue[4][20] ) );
  FDN1QM1P \Queue_reg[3][20]  ( .D(n220), .CPN(Clk_r), .Q(\Queue[3][20] ) );
  FDN1QM1P \Queue_reg[2][20]  ( .D(n252), .CPN(Clk_r), .Q(\Queue[2][20] ) );
  FDN1QM1P \Queue_reg[4][19]  ( .D(n349), .CPN(Clk_r), .Q(\Queue[4][19] ) );
  FDN1QM1P \Queue_reg[3][19]  ( .D(n221), .CPN(Clk_r), .Q(\Queue[3][19] ) );
  FDN1QM1P \Queue_reg[2][19]  ( .D(n253), .CPN(Clk_r), .Q(\Queue[2][19] ) );
  FDN1QM1P \Queue_reg[4][18]  ( .D(n350), .CPN(Clk_r), .Q(\Queue[4][18] ) );
  FDN1QM1P \Queue_reg[3][18]  ( .D(n222), .CPN(Clk_r), .Q(\Queue[3][18] ) );
  FDN1QM1P \Queue_reg[2][18]  ( .D(n254), .CPN(Clk_r), .Q(\Queue[2][18] ) );
  FDN1QM1P \Queue_reg[4][17]  ( .D(n351), .CPN(Clk_r), .Q(\Queue[4][17] ) );
  FDN1QM1P \Queue_reg[3][17]  ( .D(n223), .CPN(Clk_r), .Q(\Queue[3][17] ) );
  FDN1QM1P \Queue_reg[2][17]  ( .D(n255), .CPN(Clk_r), .Q(\Queue[2][17] ) );
  FDN1QM1P \Queue_reg[4][16]  ( .D(n352), .CPN(Clk_r), .Q(\Queue[4][16] ) );
  FDN1QM1P \Queue_reg[3][16]  ( .D(n224), .CPN(Clk_r), .Q(\Queue[3][16] ) );
  FDN1QM1P \Queue_reg[2][16]  ( .D(n256), .CPN(Clk_r), .Q(\Queue[2][16] ) );
  FDN1QM1P \Queue_reg[4][15]  ( .D(n353), .CPN(Clk_r), .Q(\Queue[4][15] ) );
  FDN1QM1P \Queue_reg[3][15]  ( .D(n225), .CPN(Clk_r), .Q(\Queue[3][15] ) );
  FDN1QM1P \Queue_reg[2][15]  ( .D(n257), .CPN(Clk_r), .Q(\Queue[2][15] ) );
  FDN1QM1P \Queue_reg[4][14]  ( .D(n354), .CPN(Clk_r), .Q(\Queue[4][14] ) );
  FDN1QM1P \Queue_reg[3][14]  ( .D(n226), .CPN(Clk_r), .Q(\Queue[3][14] ) );
  FDN1QM1P \Queue_reg[2][14]  ( .D(n258), .CPN(Clk_r), .Q(\Queue[2][14] ) );
  FDN1QM1P \Queue_reg[4][13]  ( .D(n355), .CPN(Clk_r), .Q(\Queue[4][13] ) );
  FDN1QM1P \Queue_reg[3][13]  ( .D(n227), .CPN(Clk_r), .Q(\Queue[3][13] ) );
  FDN1QM1P \Queue_reg[2][13]  ( .D(n259), .CPN(Clk_r), .Q(\Queue[2][13] ) );
  FDN1QM1P \Queue_reg[4][12]  ( .D(n356), .CPN(Clk_r), .Q(\Queue[4][12] ) );
  FDN1QM1P \Queue_reg[3][12]  ( .D(n228), .CPN(Clk_r), .Q(\Queue[3][12] ) );
  FDN1QM1P \Queue_reg[2][12]  ( .D(n260), .CPN(Clk_r), .Q(\Queue[2][12] ) );
  FDN1QM1P \Queue_reg[4][11]  ( .D(n357), .CPN(Clk_r), .Q(\Queue[4][11] ) );
  FDN1QM1P \Queue_reg[3][11]  ( .D(n229), .CPN(Clk_r), .Q(\Queue[3][11] ) );
  FDN1QM1P \Queue_reg[2][11]  ( .D(n261), .CPN(Clk_r), .Q(\Queue[2][11] ) );
  FDN1QM1P \Queue_reg[4][10]  ( .D(n358), .CPN(Clk_r), .Q(\Queue[4][10] ) );
  FDN1QM1P \Queue_reg[3][10]  ( .D(n230), .CPN(Clk_r), .Q(\Queue[3][10] ) );
  FDN1QM1P \Queue_reg[2][10]  ( .D(n262), .CPN(Clk_r), .Q(\Queue[2][10] ) );
  FDN1QM1P \Queue_reg[4][9]  ( .D(n359), .CPN(Clk_r), .Q(\Queue[4][9] ) );
  FDN1QM1P \Queue_reg[3][9]  ( .D(n231), .CPN(Clk_r), .Q(\Queue[3][9] ) );
  FDN1QM1P \Queue_reg[2][9]  ( .D(n263), .CPN(Clk_r), .Q(\Queue[2][9] ) );
  FDN1QM1P \Queue_reg[4][8]  ( .D(n360), .CPN(Clk_r), .Q(\Queue[4][8] ) );
  FDN1QM1P \Queue_reg[3][8]  ( .D(n232), .CPN(Clk_r), .Q(\Queue[3][8] ) );
  FDN1QM1P \Queue_reg[2][8]  ( .D(n264), .CPN(Clk_r), .Q(\Queue[2][8] ) );
  FDN1QM1P \Queue_reg[4][7]  ( .D(n361), .CPN(Clk_r), .Q(\Queue[4][7] ) );
  FDN1QM1P \Queue_reg[3][7]  ( .D(n233), .CPN(Clk_r), .Q(\Queue[3][7] ) );
  FDN1QM1P \Queue_reg[2][7]  ( .D(n265), .CPN(Clk_r), .Q(\Queue[2][7] ) );
  FDN1QM1P \Queue_reg[4][6]  ( .D(n362), .CPN(Clk_r), .Q(\Queue[4][6] ) );
  FDN1QM1P \Queue_reg[3][6]  ( .D(n234), .CPN(Clk_r), .Q(\Queue[3][6] ) );
  FDN1QM1P \Queue_reg[2][6]  ( .D(n266), .CPN(Clk_r), .Q(\Queue[2][6] ) );
  FDN1QM1P \Queue_reg[4][5]  ( .D(n363), .CPN(Clk_r), .Q(\Queue[4][5] ) );
  FDN1QM1P \Queue_reg[3][5]  ( .D(n235), .CPN(Clk_r), .Q(\Queue[3][5] ) );
  FDN1QM1P \Queue_reg[2][5]  ( .D(n267), .CPN(Clk_r), .Q(\Queue[2][5] ) );
  FDN1QM1P \Queue_reg[4][4]  ( .D(n364), .CPN(Clk_r), .Q(\Queue[4][4] ) );
  FDN1QM1P \Queue_reg[3][4]  ( .D(n236), .CPN(Clk_r), .Q(\Queue[3][4] ) );
  FDN1QM1P \Queue_reg[2][4]  ( .D(n268), .CPN(Clk_r), .Q(\Queue[2][4] ) );
  FDN1QM1P \Queue_reg[4][3]  ( .D(n365), .CPN(Clk_r), .Q(\Queue[4][3] ) );
  FDN1QM1P \Queue_reg[3][3]  ( .D(n237), .CPN(Clk_r), .Q(\Queue[3][3] ) );
  FDN1QM1P \Queue_reg[2][3]  ( .D(n269), .CPN(Clk_r), .Q(\Queue[2][3] ) );
  FDN1QM1P \Queue_reg[4][2]  ( .D(n366), .CPN(Clk_r), .Q(\Queue[4][2] ) );
  FDN1QM1P \Queue_reg[3][2]  ( .D(n238), .CPN(Clk_r), .Q(\Queue[3][2] ) );
  FDN1QM1P \Queue_reg[2][2]  ( .D(n270), .CPN(Clk_r), .Q(\Queue[2][2] ) );
  FDN1QM1P \Queue_reg[4][1]  ( .D(n367), .CPN(Clk_r), .Q(\Queue[4][1] ) );
  FDN1QM1P \Queue_reg[3][1]  ( .D(n239), .CPN(Clk_r), .Q(\Queue[3][1] ) );
  FDN1QM1P \Queue_reg[2][1]  ( .D(n271), .CPN(Clk_r), .Q(\Queue[2][1] ) );
  FDN1QM1P \Queue_reg[4][0]  ( .D(n368), .CPN(Clk_r), .Q(\Queue[4][0] ) );
  FDN1QM1P \Queue_reg[3][0]  ( .D(n240), .CPN(Clk_r), .Q(\Queue[3][0] ) );
  FDN1QM1P \Queue_reg[2][0]  ( .D(n272), .CPN(Clk_r), .Q(\Queue[2][0] ) );
  FDN1QM1P \Queue_reg[4][31]  ( .D(n369), .CPN(Clk_r), .Q(\Queue[4][31] ) );
  FDN1QM1P \Queue_reg[3][31]  ( .D(n209), .CPN(Clk_r), .Q(\Queue[3][31] ) );
  FDN1QM1P \Queue_reg[2][31]  ( .D(n241), .CPN(Clk_r), .Q(\Queue[2][31] ) );
  FDN2QM1P Full_reg ( .D(n337), .CPN(Clk_r), .CD(Rst_n), .Q(Full) );
  FDN1QM1P \Queue_reg[1][31]  ( .D(n305), .CPN(Clk_r), .Q(\Queue[1][31] ) );
  FDN1QM1P \Queue_reg[0][31]  ( .D(n273), .CPN(Clk_r), .Q(Packet_Out[31]) );
  FDN1QM1P \Queue_reg[1][30]  ( .D(n306), .CPN(Clk_r), .Q(\Queue[1][30] ) );
  FDN1QM1P \Queue_reg[0][30]  ( .D(n274), .CPN(Clk_r), .Q(Packet_Out[30]) );
  FDN1QM1P \Queue_reg[1][29]  ( .D(n307), .CPN(Clk_r), .Q(\Queue[1][29] ) );
  FDN1QM1P \Queue_reg[0][29]  ( .D(n275), .CPN(Clk_r), .Q(Packet_Out[29]) );
  FDN1QM1P \Queue_reg[1][28]  ( .D(n308), .CPN(Clk_r), .Q(\Queue[1][28] ) );
  FDN1QM1P \Queue_reg[0][28]  ( .D(n276), .CPN(Clk_r), .Q(Packet_Out[28]) );
  FDN1QM1P \Queue_reg[1][27]  ( .D(n309), .CPN(Clk_r), .Q(\Queue[1][27] ) );
  FDN1QM1P \Queue_reg[0][27]  ( .D(n277), .CPN(Clk_r), .Q(Packet_Out[27]) );
  FDN1QM1P \Queue_reg[1][26]  ( .D(n310), .CPN(Clk_r), .Q(\Queue[1][26] ) );
  FDN1QM1P \Queue_reg[0][26]  ( .D(n278), .CPN(Clk_r), .Q(Packet_Out[26]) );
  FDN1QM1P \Queue_reg[1][25]  ( .D(n311), .CPN(Clk_r), .Q(\Queue[1][25] ) );
  FDN1QM1P \Queue_reg[0][25]  ( .D(n279), .CPN(Clk_r), .Q(Packet_Out[25]) );
  FDN1QM1P \Queue_reg[1][24]  ( .D(n312), .CPN(Clk_r), .Q(\Queue[1][24] ) );
  FDN1QM1P \Queue_reg[0][24]  ( .D(n280), .CPN(Clk_r), .Q(Packet_Out[24]) );
  FDN1QM1P \Queue_reg[1][23]  ( .D(n313), .CPN(Clk_r), .Q(\Queue[1][23] ) );
  FDN1QM1P \Queue_reg[0][23]  ( .D(n281), .CPN(Clk_r), .Q(Packet_Out[23]) );
  FDN1QM1P \Queue_reg[1][22]  ( .D(n314), .CPN(Clk_r), .Q(\Queue[1][22] ) );
  FDN1QM1P \Queue_reg[0][22]  ( .D(n282), .CPN(Clk_r), .Q(Packet_Out[22]) );
  FDN1QM1P \Queue_reg[1][21]  ( .D(n315), .CPN(Clk_r), .Q(\Queue[1][21] ) );
  FDN1QM1P \Queue_reg[0][21]  ( .D(n283), .CPN(Clk_r), .Q(Packet_Out[21]) );
  FDN1QM1P \Queue_reg[1][20]  ( .D(n316), .CPN(Clk_r), .Q(\Queue[1][20] ) );
  FDN1QM1P \Queue_reg[0][20]  ( .D(n284), .CPN(Clk_r), .Q(Packet_Out[20]) );
  FDN1QM1P \Queue_reg[1][19]  ( .D(n317), .CPN(Clk_r), .Q(\Queue[1][19] ) );
  FDN1QM1P \Queue_reg[0][19]  ( .D(n285), .CPN(Clk_r), .Q(Packet_Out[19]) );
  FDN1QM1P \Queue_reg[1][18]  ( .D(n318), .CPN(Clk_r), .Q(\Queue[1][18] ) );
  FDN1QM1P \Queue_reg[0][18]  ( .D(n286), .CPN(Clk_r), .Q(Packet_Out[18]) );
  FDN1QM1P \Queue_reg[1][17]  ( .D(n319), .CPN(Clk_r), .Q(\Queue[1][17] ) );
  FDN1QM1P \Queue_reg[0][17]  ( .D(n287), .CPN(Clk_r), .Q(Packet_Out[17]) );
  FDN1QM1P \Queue_reg[1][16]  ( .D(n320), .CPN(Clk_r), .Q(\Queue[1][16] ) );
  FDN1QM1P \Queue_reg[0][16]  ( .D(n288), .CPN(Clk_r), .Q(Packet_Out[16]) );
  FDN1QM1P \Queue_reg[1][15]  ( .D(n321), .CPN(Clk_r), .Q(\Queue[1][15] ) );
  FDN1QM1P \Queue_reg[0][15]  ( .D(n289), .CPN(Clk_r), .Q(Packet_Out[15]) );
  FDN1QM1P \Queue_reg[1][14]  ( .D(n322), .CPN(Clk_r), .Q(\Queue[1][14] ) );
  FDN1QM1P \Queue_reg[0][14]  ( .D(n290), .CPN(Clk_r), .Q(Packet_Out[14]) );
  FDN1QM1P \Queue_reg[1][13]  ( .D(n323), .CPN(Clk_r), .Q(\Queue[1][13] ) );
  FDN1QM1P \Queue_reg[0][13]  ( .D(n291), .CPN(Clk_r), .Q(Packet_Out[13]) );
  FDN1QM1P \Queue_reg[1][12]  ( .D(n324), .CPN(Clk_r), .Q(\Queue[1][12] ) );
  FDN1QM1P \Queue_reg[0][12]  ( .D(n292), .CPN(Clk_r), .Q(Packet_Out[12]) );
  FDN1QM1P \Queue_reg[1][11]  ( .D(n325), .CPN(Clk_r), .Q(\Queue[1][11] ) );
  FDN1QM1P \Queue_reg[0][11]  ( .D(n293), .CPN(Clk_r), .Q(Packet_Out[11]) );
  FDN1QM1P \Queue_reg[1][10]  ( .D(n326), .CPN(Clk_r), .Q(\Queue[1][10] ) );
  FDN1QM1P \Queue_reg[0][10]  ( .D(n294), .CPN(Clk_r), .Q(Packet_Out[10]) );
  FDN1QM1P \Queue_reg[1][9]  ( .D(n327), .CPN(Clk_r), .Q(\Queue[1][9] ) );
  FDN1QM1P \Queue_reg[0][9]  ( .D(n295), .CPN(Clk_r), .Q(Packet_Out[9]) );
  FDN1QM1P \Queue_reg[1][8]  ( .D(n328), .CPN(Clk_r), .Q(\Queue[1][8] ) );
  FDN1QM1P \Queue_reg[0][8]  ( .D(n296), .CPN(Clk_r), .Q(Packet_Out[8]) );
  FDN1QM1P \Queue_reg[1][7]  ( .D(n329), .CPN(Clk_r), .Q(\Queue[1][7] ) );
  FDN1QM1P \Queue_reg[0][7]  ( .D(n297), .CPN(Clk_r), .Q(Packet_Out[7]) );
  FDN1QM1P \Queue_reg[1][6]  ( .D(n330), .CPN(Clk_r), .Q(\Queue[1][6] ) );
  FDN1QM1P \Queue_reg[0][6]  ( .D(n298), .CPN(Clk_r), .Q(Packet_Out[6]) );
  FDN1QM1P \Queue_reg[1][5]  ( .D(n331), .CPN(Clk_r), .Q(\Queue[1][5] ) );
  FDN1QM1P \Queue_reg[0][5]  ( .D(n299), .CPN(Clk_r), .Q(Packet_Out[5]) );
  FDN1QM1P \Queue_reg[1][4]  ( .D(n332), .CPN(Clk_r), .Q(\Queue[1][4] ) );
  FDN1QM1P \Queue_reg[0][4]  ( .D(n300), .CPN(Clk_r), .Q(Packet_Out[4]) );
  FDN1QM1P \Queue_reg[1][3]  ( .D(n333), .CPN(Clk_r), .Q(\Queue[1][3] ) );
  FDN1QM1P \Queue_reg[0][3]  ( .D(n301), .CPN(Clk_r), .Q(Packet_Out[3]) );
  FDN1QM1P \Queue_reg[1][2]  ( .D(n334), .CPN(Clk_r), .Q(\Queue[1][2] ) );
  FDN1QM1P \Queue_reg[0][2]  ( .D(n302), .CPN(Clk_r), .Q(Packet_Out[2]) );
  FDN1QM1P \Queue_reg[1][1]  ( .D(n335), .CPN(Clk_r), .Q(\Queue[1][1] ) );
  FDN1QM1P \Queue_reg[0][1]  ( .D(n303), .CPN(Clk_r), .Q(Packet_Out[1]) );
  FDN1QM1P \Queue_reg[1][0]  ( .D(n336), .CPN(Clk_r), .Q(\Queue[1][0] ) );
  FDN1QM1P \Queue_reg[0][0]  ( .D(n304), .CPN(Clk_r), .Q(Packet_Out[0]) );
  FDN2QM1P Empty_reg ( .D(n1), .CPN(Clk_r), .CD(Rst_n), .Q(n2) );
  NR3M1P U3 ( .A(Count[0]), .B(Count[2]), .C(n22), .Z(n100) );
  N1M1P U4 ( .A(Read_Ack), .Z(n137) );
  BUFM2P U5 ( .A(n95), .Z(n3) );
  BUFM2P U6 ( .A(n132), .Z(n5) );
  BUFM2P U7 ( .A(n205), .Z(n4) );
  NR3M1P U8 ( .A(n23), .B(Count[2]), .C(Count[1]), .Z(n376) );
  NR3M1P U9 ( .A(Count[2]), .B(n23), .C(n22), .Z(n140) );
  OAI21M2P U10 ( .A(n61), .B(n60), .C(n141), .Z(n62) );
  AOI21M6P U11 ( .A(n6), .B(n100), .C(n141), .Z(n57) );
  BUFM1P U12 ( .A(n57), .Z(n9) );
  OAI211M4P U13 ( .A(n140), .B(n137), .C(n6), .D(n98), .Z(n135) );
  OAI211M4P U14 ( .A(n142), .B(n137), .C(n6), .D(n136), .Z(n208) );
  BUFM2P U15 ( .A(n97), .Z(n12) );
  NR2FM3P U16 ( .A(n61), .B(n21), .Z(n20) );
  OAI211M4P U17 ( .A(n100), .B(n139), .C(Rst_n), .D(n138), .Z(n133) );
  OAI211M4P U18 ( .A(n140), .B(n139), .C(Rst_n), .D(n138), .Z(n206) );
  OAI21M2P U19 ( .A(n6), .B(Read_Ack), .C(n24), .Z(n56) );
  NR3M1P U20 ( .A(Count[0]), .B(Count[1]), .C(n19), .Z(n142) );
  N1M2P U21 ( .A(n6), .Z(n99) );
  N1M1P U22 ( .A(Count[1]), .Z(n22) );
  N1M1P U23 ( .A(Count[2]), .Z(n19) );
  N1M1P U24 ( .A(Count[0]), .Z(n23) );
  ND2M2P U25 ( .A(n18), .B(Rst_n), .Z(n61) );
  ND2M2P U26 ( .A(Read_Ack), .B(Rst_n), .Z(n141) );
  OAI211M2P U27 ( .A(n100), .B(n137), .C(n6), .D(n24), .Z(n59) );
  NR2FM2P U28 ( .A(Read_Ack), .B(n99), .Z(n18) );
  N1M1P U29 ( .A(Packet_In[29]), .Z(n202) );
  N1M1P U30 ( .A(Packet_In[0]), .Z(n144) );
  N1M1P U31 ( .A(Packet_In[8]), .Z(n160) );
  N1M1P U32 ( .A(Packet_In[3]), .Z(n150) );
  N1M1P U33 ( .A(Packet_In[4]), .Z(n152) );
  N1M1P U34 ( .A(Packet_In[5]), .Z(n154) );
  N1M1P U35 ( .A(Packet_In[6]), .Z(n156) );
  N1M1P U36 ( .A(Packet_In[7]), .Z(n158) );
  N1M1P U37 ( .A(Packet_In[2]), .Z(n148) );
  N1M1P U38 ( .A(Packet_In[1]), .Z(n146) );
  N1M1P U39 ( .A(Packet_In[26]), .Z(n196) );
  N1M1P U40 ( .A(Packet_In[25]), .Z(n194) );
  N1M1P U41 ( .A(Packet_In[31]), .Z(n373) );
  N1M1P U42 ( .A(Packet_In[30]), .Z(n204) );
  N1M1P U43 ( .A(Packet_In[28]), .Z(n200) );
  N1M1P U44 ( .A(Packet_In[27]), .Z(n198) );
  N1M1P U45 ( .A(Packet_In[20]), .Z(n184) );
  N1M1P U46 ( .A(Packet_In[17]), .Z(n178) );
  N1M1P U47 ( .A(Packet_In[16]), .Z(n176) );
  N1M1P U48 ( .A(Packet_In[15]), .Z(n174) );
  N1M1P U49 ( .A(Packet_In[19]), .Z(n182) );
  N1M1P U50 ( .A(Packet_In[13]), .Z(n170) );
  N1M1P U51 ( .A(Packet_In[23]), .Z(n190) );
  N1M1P U52 ( .A(Packet_In[12]), .Z(n168) );
  N1M1P U53 ( .A(Packet_In[18]), .Z(n180) );
  N1M1P U54 ( .A(Packet_In[14]), .Z(n172) );
  N1M1P U55 ( .A(Packet_In[21]), .Z(n186) );
  N1M1P U56 ( .A(Packet_In[9]), .Z(n162) );
  N1M1P U57 ( .A(Packet_In[22]), .Z(n188) );
  N1M1P U58 ( .A(Packet_In[10]), .Z(n164) );
  N1M1P U59 ( .A(Packet_In[24]), .Z(n192) );
  N1M1P U60 ( .A(Packet_In[11]), .Z(n166) );
  N1M2P U61 ( .A(n62), .Z(n94) );
  OAI211M1P U62 ( .A(n376), .B(n137), .C(n6), .D(n62), .Z(n97) );
  BUFM2P U63 ( .A(n59), .Z(n11) );
  BUFM2P U64 ( .A(n56), .Z(n8) );
  BUFM2P U65 ( .A(n59), .Z(n10) );
  BUFM2P U66 ( .A(n56), .Z(n7) );
  N1M2P U67 ( .A(n18), .Z(n139) );
  BUFM6P U68 ( .A(Write_Ack), .Z(n6) );
  AOI22M1P U69 ( .A(\Queue[2][1] ), .B(n133), .C(n5), .D(\Queue[3][1] ), .Z(
        n102) );
  NR2M1P U70 ( .A(n137), .B(n6), .Z(n375) );
  NR2M1P U71 ( .A(n18), .B(n375), .Z(n374) );
  AOI22CDNM1P U72 ( .A(n374), .B(n23), .C(n374), .D(n23), .Z(n372) );
  N1M1P U73 ( .A(n375), .Z(n17) );
  AOI22M1P U74 ( .A(Count[0]), .B(n139), .C(n17), .D(n23), .Z(n14) );
  AOI22CDNM1P U75 ( .A(Count[1]), .B(n14), .C(n14), .D(Count[1]), .Z(n371) );
  ND3M1P U76 ( .A(n23), .B(n19), .C(n22), .Z(n60) );
  ND2M1P U77 ( .A(Count[1]), .B(Read_Ack), .Z(n13) );
  OAI211M1P U78 ( .A(Count[1]), .B(n139), .C(n14), .D(n13), .Z(n15) );
  AOI22M1P U79 ( .A(n18), .B(n140), .C(Count[2]), .D(n15), .Z(n16) );
  OAI21M1P U80 ( .A(n60), .B(n17), .C(n16), .Z(n370) );
  N1M1P U81 ( .A(n142), .Z(n21) );
  AOI22CDNM1P U82 ( .A(n20), .B(n373), .C(\Queue[4][31] ), .D(n20), .Z(n369)
         );
  AOI22CDNM1P U83 ( .A(n20), .B(n144), .C(\Queue[4][0] ), .D(n20), .Z(n368) );
  AOI22CDNM1P U84 ( .A(n20), .B(n146), .C(\Queue[4][1] ), .D(n20), .Z(n367) );
  AOI22CDNM1P U85 ( .A(n20), .B(n148), .C(\Queue[4][2] ), .D(n20), .Z(n366) );
  AOI22CDNM1P U86 ( .A(n20), .B(n150), .C(\Queue[4][3] ), .D(n20), .Z(n365) );
  AOI22CDNM1P U87 ( .A(n20), .B(n152), .C(\Queue[4][4] ), .D(n20), .Z(n364) );
  AOI22CDNM1P U88 ( .A(n20), .B(n154), .C(\Queue[4][5] ), .D(n20), .Z(n363) );
  AOI22CDNM1P U89 ( .A(n20), .B(n156), .C(\Queue[4][6] ), .D(n20), .Z(n362) );
  AOI22CDNM1P U90 ( .A(n20), .B(n158), .C(\Queue[4][7] ), .D(n20), .Z(n361) );
  AOI22CDNM1P U91 ( .A(n20), .B(n160), .C(\Queue[4][8] ), .D(n20), .Z(n360) );
  AOI22CDNM1P U92 ( .A(n20), .B(n162), .C(\Queue[4][9] ), .D(n20), .Z(n359) );
  AOI22CDNM1P U93 ( .A(n20), .B(n164), .C(\Queue[4][10] ), .D(n20), .Z(n358)
         );
  AOI22CDNM1P U94 ( .A(n20), .B(n166), .C(\Queue[4][11] ), .D(n20), .Z(n357)
         );
  AOI22CDNM1P U95 ( .A(n20), .B(n168), .C(\Queue[4][12] ), .D(n20), .Z(n356)
         );
  AOI22CDNM1P U96 ( .A(n20), .B(n170), .C(\Queue[4][13] ), .D(n20), .Z(n355)
         );
  AOI22CDNM1P U97 ( .A(n20), .B(n172), .C(\Queue[4][14] ), .D(n20), .Z(n354)
         );
  AOI22CDNM1P U98 ( .A(n20), .B(n174), .C(\Queue[4][15] ), .D(n20), .Z(n353)
         );
  AOI22CDNM1P U99 ( .A(n20), .B(n176), .C(\Queue[4][16] ), .D(n20), .Z(n352)
         );
  AOI22CDNM1P U100 ( .A(n20), .B(n178), .C(\Queue[4][17] ), .D(n20), .Z(n351)
         );
  AOI22CDNM1P U101 ( .A(n20), .B(n180), .C(\Queue[4][18] ), .D(n20), .Z(n350)
         );
  AOI22CDNM1P U102 ( .A(n20), .B(n182), .C(\Queue[4][19] ), .D(n20), .Z(n349)
         );
  AOI22CDNM1P U103 ( .A(n20), .B(n184), .C(\Queue[4][20] ), .D(n20), .Z(n348)
         );
  AOI22CDNM1P U104 ( .A(n20), .B(n186), .C(\Queue[4][21] ), .D(n20), .Z(n347)
         );
  AOI22CDNM1P U105 ( .A(n20), .B(n188), .C(\Queue[4][22] ), .D(n20), .Z(n346)
         );
  AOI22CDNM1P U106 ( .A(n20), .B(n190), .C(\Queue[4][23] ), .D(n20), .Z(n345)
         );
  AOI22CDNM1P U107 ( .A(n20), .B(n192), .C(\Queue[4][24] ), .D(n20), .Z(n344)
         );
  AOI22CDNM1P U108 ( .A(n20), .B(n194), .C(\Queue[4][25] ), .D(n20), .Z(n343)
         );
  AOI22CDNM1P U109 ( .A(n20), .B(n196), .C(\Queue[4][26] ), .D(n20), .Z(n342)
         );
  AOI22CDNM1P U110 ( .A(n20), .B(n198), .C(\Queue[4][27] ), .D(n20), .Z(n341)
         );
  AOI22CDNM1P U111 ( .A(n20), .B(n200), .C(\Queue[4][28] ), .D(n20), .Z(n340)
         );
  AOI22CDNM1P U112 ( .A(n20), .B(n202), .C(\Queue[4][29] ), .D(n20), .Z(n339)
         );
  AOI22CDNM1P U113 ( .A(n20), .B(n204), .C(\Queue[4][30] ), .D(n20), .Z(n338)
         );
  OAI22CDNM1P U114 ( .A(n139), .B(n21), .C(n374), .D(Full), .Z(n337) );
  OA21M1P U115 ( .A(n139), .B(n376), .C(Rst_n), .Z(n24) );
  AOI22M1P U116 ( .A(\Queue[2][0] ), .B(n57), .C(\Queue[1][0] ), .D(n56), .Z(
        n25) );
  OAI21M1P U117 ( .A(n144), .B(n59), .C(n25), .Z(n336) );
  AOI22M1P U118 ( .A(n9), .B(\Queue[2][1] ), .C(\Queue[1][1] ), .D(n7), .Z(n26) );
  OAI21M1P U119 ( .A(n59), .B(n146), .C(n26), .Z(n335) );
  AOI22M1P U120 ( .A(n57), .B(\Queue[2][2] ), .C(\Queue[1][2] ), .D(n56), .Z(
        n27) );
  OAI21M1P U121 ( .A(n10), .B(n148), .C(n27), .Z(n334) );
  AOI22M1P U122 ( .A(n57), .B(\Queue[2][3] ), .C(\Queue[1][3] ), .D(n56), .Z(
        n28) );
  OAI21M1P U123 ( .A(n11), .B(n150), .C(n28), .Z(n333) );
  AOI22M1P U124 ( .A(n57), .B(\Queue[2][4] ), .C(\Queue[1][4] ), .D(n56), .Z(
        n29) );
  OAI21M1P U125 ( .A(n10), .B(n152), .C(n29), .Z(n332) );
  AOI22M1P U126 ( .A(n57), .B(\Queue[2][5] ), .C(\Queue[1][5] ), .D(n56), .Z(
        n30) );
  OAI21M1P U127 ( .A(n11), .B(n154), .C(n30), .Z(n331) );
  AOI22M1P U128 ( .A(n9), .B(\Queue[2][6] ), .C(\Queue[1][6] ), .D(n56), .Z(
        n31) );
  OAI21M1P U129 ( .A(n59), .B(n156), .C(n31), .Z(n330) );
  AOI22M1P U130 ( .A(n57), .B(\Queue[2][7] ), .C(\Queue[1][7] ), .D(n56), .Z(
        n32) );
  OAI21M1P U131 ( .A(n59), .B(n158), .C(n32), .Z(n329) );
  AOI22M1P U132 ( .A(n57), .B(\Queue[2][8] ), .C(\Queue[1][8] ), .D(n56), .Z(
        n33) );
  OAI21M1P U133 ( .A(n59), .B(n160), .C(n33), .Z(n328) );
  AOI22M1P U134 ( .A(n57), .B(\Queue[2][9] ), .C(\Queue[1][9] ), .D(n7), .Z(
        n34) );
  OAI21M1P U135 ( .A(n59), .B(n162), .C(n34), .Z(n327) );
  AOI22M1P U136 ( .A(n57), .B(\Queue[2][10] ), .C(\Queue[1][10] ), .D(n7), .Z(
        n35) );
  OAI21M1P U137 ( .A(n59), .B(n164), .C(n35), .Z(n326) );
  AOI22M1P U138 ( .A(n57), .B(\Queue[2][11] ), .C(\Queue[1][11] ), .D(n7), .Z(
        n36) );
  OAI21M1P U139 ( .A(n59), .B(n166), .C(n36), .Z(n325) );
  AOI22M1P U140 ( .A(n9), .B(\Queue[2][12] ), .C(\Queue[1][12] ), .D(n7), .Z(
        n37) );
  OAI21M1P U141 ( .A(n11), .B(n168), .C(n37), .Z(n324) );
  AOI22M1P U142 ( .A(n9), .B(\Queue[2][13] ), .C(\Queue[1][13] ), .D(n7), .Z(
        n38) );
  OAI21M1P U143 ( .A(n11), .B(n170), .C(n38), .Z(n323) );
  AOI22M1P U144 ( .A(n9), .B(\Queue[2][14] ), .C(\Queue[1][14] ), .D(n7), .Z(
        n39) );
  OAI21M1P U145 ( .A(n11), .B(n172), .C(n39), .Z(n322) );
  AOI22M1P U146 ( .A(n9), .B(\Queue[2][15] ), .C(\Queue[1][15] ), .D(n7), .Z(
        n40) );
  OAI21M1P U147 ( .A(n11), .B(n174), .C(n40), .Z(n321) );
  AOI22M1P U148 ( .A(n9), .B(\Queue[2][16] ), .C(\Queue[1][16] ), .D(n7), .Z(
        n41) );
  OAI21M1P U149 ( .A(n11), .B(n176), .C(n41), .Z(n320) );
  AOI22M1P U150 ( .A(n9), .B(\Queue[2][17] ), .C(\Queue[1][17] ), .D(n7), .Z(
        n42) );
  OAI21M1P U151 ( .A(n11), .B(n178), .C(n42), .Z(n319) );
  AOI22M1P U152 ( .A(n9), .B(\Queue[2][18] ), .C(\Queue[1][18] ), .D(n8), .Z(
        n43) );
  OAI21M1P U153 ( .A(n11), .B(n180), .C(n43), .Z(n318) );
  AOI22M1P U154 ( .A(n9), .B(\Queue[2][19] ), .C(\Queue[1][19] ), .D(n8), .Z(
        n44) );
  OAI21M1P U155 ( .A(n11), .B(n182), .C(n44), .Z(n317) );
  AOI22M1P U156 ( .A(n9), .B(\Queue[2][20] ), .C(\Queue[1][20] ), .D(n8), .Z(
        n45) );
  OAI21M1P U157 ( .A(n11), .B(n184), .C(n45), .Z(n316) );
  AOI22M1P U158 ( .A(n9), .B(\Queue[2][21] ), .C(\Queue[1][21] ), .D(n8), .Z(
        n46) );
  OAI21M1P U159 ( .A(n11), .B(n186), .C(n46), .Z(n315) );
  AOI22M1P U160 ( .A(n57), .B(\Queue[2][22] ), .C(\Queue[1][22] ), .D(n8), .Z(
        n47) );
  OAI21M1P U161 ( .A(n10), .B(n188), .C(n47), .Z(n314) );
  AOI22M1P U162 ( .A(n9), .B(\Queue[2][23] ), .C(\Queue[1][23] ), .D(n8), .Z(
        n48) );
  OAI21M1P U163 ( .A(n10), .B(n190), .C(n48), .Z(n313) );
  AOI22M1P U164 ( .A(n57), .B(\Queue[2][24] ), .C(\Queue[1][24] ), .D(n8), .Z(
        n49) );
  OAI21M1P U165 ( .A(n10), .B(n192), .C(n49), .Z(n312) );
  AOI22M1P U166 ( .A(n57), .B(\Queue[2][25] ), .C(\Queue[1][25] ), .D(n8), .Z(
        n50) );
  OAI21M1P U167 ( .A(n10), .B(n194), .C(n50), .Z(n311) );
  AOI22M1P U168 ( .A(n57), .B(\Queue[2][26] ), .C(\Queue[1][26] ), .D(n8), .Z(
        n51) );
  OAI21M1P U169 ( .A(n10), .B(n196), .C(n51), .Z(n310) );
  AOI22M1P U170 ( .A(n57), .B(\Queue[2][27] ), .C(\Queue[1][27] ), .D(n7), .Z(
        n52) );
  OAI21M1P U171 ( .A(n10), .B(n198), .C(n52), .Z(n309) );
  AOI22M1P U172 ( .A(n57), .B(\Queue[2][28] ), .C(\Queue[1][28] ), .D(n8), .Z(
        n53) );
  OAI21M1P U173 ( .A(n10), .B(n200), .C(n53), .Z(n308) );
  AOI22M1P U174 ( .A(n57), .B(\Queue[2][29] ), .C(\Queue[1][29] ), .D(n8), .Z(
        n54) );
  OAI21M1P U175 ( .A(n10), .B(n202), .C(n54), .Z(n307) );
  AOI22M1P U176 ( .A(n57), .B(\Queue[2][30] ), .C(\Queue[1][30] ), .D(n7), .Z(
        n55) );
  OAI21M1P U177 ( .A(n10), .B(n204), .C(n55), .Z(n306) );
  AOI22M1P U178 ( .A(n57), .B(\Queue[2][31] ), .C(\Queue[1][31] ), .D(n8), .Z(
        n58) );
  OAI21M1P U179 ( .A(n10), .B(n373), .C(n58), .Z(n305) );
  AOI21M1P U180 ( .A(n6), .B(n376), .C(n141), .Z(n95) );
  AOI22M1P U181 ( .A(\Queue[1][0] ), .B(n3), .C(n94), .D(Packet_Out[0]), .Z(
        n63) );
  OAI21M1P U182 ( .A(n144), .B(n12), .C(n63), .Z(n304) );
  AOI22M1P U183 ( .A(\Queue[1][1] ), .B(n3), .C(n94), .D(Packet_Out[1]), .Z(
        n64) );
  OAI21M1P U184 ( .A(n146), .B(n12), .C(n64), .Z(n303) );
  AOI22M1P U185 ( .A(\Queue[1][2] ), .B(n3), .C(n94), .D(Packet_Out[2]), .Z(
        n65) );
  OAI21M1P U186 ( .A(n148), .B(n12), .C(n65), .Z(n302) );
  AOI22M1P U187 ( .A(\Queue[1][3] ), .B(n3), .C(n94), .D(Packet_Out[3]), .Z(
        n66) );
  OAI21M1P U188 ( .A(n150), .B(n12), .C(n66), .Z(n301) );
  AOI22M1P U189 ( .A(\Queue[1][4] ), .B(n3), .C(n94), .D(Packet_Out[4]), .Z(
        n67) );
  OAI21M1P U190 ( .A(n152), .B(n12), .C(n67), .Z(n300) );
  AOI22M1P U191 ( .A(\Queue[1][5] ), .B(n3), .C(n94), .D(Packet_Out[5]), .Z(
        n68) );
  OAI21M1P U192 ( .A(n154), .B(n12), .C(n68), .Z(n299) );
  AOI22M1P U193 ( .A(\Queue[1][6] ), .B(n3), .C(n94), .D(Packet_Out[6]), .Z(
        n69) );
  OAI21M1P U194 ( .A(n156), .B(n12), .C(n69), .Z(n298) );
  AOI22M1P U195 ( .A(\Queue[1][7] ), .B(n3), .C(n94), .D(Packet_Out[7]), .Z(
        n70) );
  OAI21M1P U196 ( .A(n158), .B(n12), .C(n70), .Z(n297) );
  AOI22M1P U197 ( .A(\Queue[1][8] ), .B(n3), .C(n94), .D(Packet_Out[8]), .Z(
        n71) );
  OAI21M1P U198 ( .A(n160), .B(n12), .C(n71), .Z(n296) );
  AOI22M1P U199 ( .A(\Queue[1][9] ), .B(n3), .C(n94), .D(Packet_Out[9]), .Z(
        n72) );
  OAI21M1P U200 ( .A(n162), .B(n12), .C(n72), .Z(n295) );
  AOI22M1P U201 ( .A(\Queue[1][10] ), .B(n3), .C(n94), .D(Packet_Out[10]), .Z(
        n73) );
  OAI21M1P U202 ( .A(n164), .B(n12), .C(n73), .Z(n294) );
  AOI22M1P U203 ( .A(\Queue[1][11] ), .B(n3), .C(n94), .D(Packet_Out[11]), .Z(
        n74) );
  OAI21M1P U204 ( .A(n166), .B(n12), .C(n74), .Z(n293) );
  AOI22M1P U205 ( .A(\Queue[1][12] ), .B(n3), .C(n94), .D(Packet_Out[12]), .Z(
        n75) );
  OAI21M1P U206 ( .A(n168), .B(n12), .C(n75), .Z(n292) );
  AOI22M1P U207 ( .A(\Queue[1][13] ), .B(n3), .C(n94), .D(Packet_Out[13]), .Z(
        n76) );
  OAI21M1P U208 ( .A(n170), .B(n12), .C(n76), .Z(n291) );
  AOI22M1P U209 ( .A(\Queue[1][14] ), .B(n3), .C(n94), .D(Packet_Out[14]), .Z(
        n77) );
  OAI21M1P U210 ( .A(n172), .B(n12), .C(n77), .Z(n290) );
  AOI22M1P U211 ( .A(\Queue[1][15] ), .B(n3), .C(n94), .D(Packet_Out[15]), .Z(
        n78) );
  OAI21M1P U212 ( .A(n174), .B(n12), .C(n78), .Z(n289) );
  AOI22M1P U213 ( .A(\Queue[1][16] ), .B(n3), .C(n94), .D(Packet_Out[16]), .Z(
        n79) );
  OAI21M1P U214 ( .A(n176), .B(n12), .C(n79), .Z(n288) );
  AOI22M1P U215 ( .A(\Queue[1][17] ), .B(n3), .C(n94), .D(Packet_Out[17]), .Z(
        n80) );
  OAI21M1P U216 ( .A(n178), .B(n12), .C(n80), .Z(n287) );
  AOI22M1P U217 ( .A(\Queue[1][18] ), .B(n3), .C(n94), .D(Packet_Out[18]), .Z(
        n81) );
  OAI21M1P U218 ( .A(n180), .B(n12), .C(n81), .Z(n286) );
  AOI22M1P U219 ( .A(\Queue[1][19] ), .B(n3), .C(n94), .D(Packet_Out[19]), .Z(
        n82) );
  OAI21M1P U220 ( .A(n182), .B(n12), .C(n82), .Z(n285) );
  AOI22M1P U221 ( .A(\Queue[1][20] ), .B(n3), .C(n94), .D(Packet_Out[20]), .Z(
        n83) );
  OAI21M1P U222 ( .A(n184), .B(n97), .C(n83), .Z(n284) );
  AOI22M1P U223 ( .A(\Queue[1][21] ), .B(n3), .C(n94), .D(Packet_Out[21]), .Z(
        n84) );
  OAI21M1P U224 ( .A(n186), .B(n97), .C(n84), .Z(n283) );
  AOI22M1P U225 ( .A(\Queue[1][22] ), .B(n3), .C(n94), .D(Packet_Out[22]), .Z(
        n85) );
  OAI21M1P U226 ( .A(n188), .B(n12), .C(n85), .Z(n282) );
  AOI22M1P U227 ( .A(\Queue[1][23] ), .B(n3), .C(n94), .D(Packet_Out[23]), .Z(
        n86) );
  OAI21M1P U228 ( .A(n190), .B(n12), .C(n86), .Z(n281) );
  AOI22M1P U229 ( .A(\Queue[1][24] ), .B(n3), .C(n94), .D(Packet_Out[24]), .Z(
        n87) );
  OAI21M1P U230 ( .A(n192), .B(n12), .C(n87), .Z(n280) );
  AOI22M1P U231 ( .A(\Queue[1][25] ), .B(n3), .C(n94), .D(Packet_Out[25]), .Z(
        n88) );
  OAI21M1P U232 ( .A(n194), .B(n12), .C(n88), .Z(n279) );
  AOI22M1P U233 ( .A(\Queue[1][26] ), .B(n3), .C(n94), .D(Packet_Out[26]), .Z(
        n89) );
  OAI21M1P U234 ( .A(n196), .B(n12), .C(n89), .Z(n278) );
  AOI22M1P U235 ( .A(\Queue[1][27] ), .B(n3), .C(n94), .D(Packet_Out[27]), .Z(
        n90) );
  OAI21M1P U236 ( .A(n198), .B(n12), .C(n90), .Z(n277) );
  AOI22M1P U237 ( .A(\Queue[1][28] ), .B(n3), .C(n94), .D(Packet_Out[28]), .Z(
        n91) );
  OAI21M1P U238 ( .A(n200), .B(n12), .C(n91), .Z(n276) );
  AOI22M1P U239 ( .A(\Queue[1][29] ), .B(n3), .C(n94), .D(Packet_Out[29]), .Z(
        n92) );
  OAI21M1P U240 ( .A(n202), .B(n12), .C(n92), .Z(n275) );
  AOI22M1P U241 ( .A(\Queue[1][30] ), .B(n95), .C(n94), .D(Packet_Out[30]), 
        .Z(n93) );
  OAI21M1P U242 ( .A(n204), .B(n12), .C(n93), .Z(n274) );
  AOI22M1P U243 ( .A(\Queue[1][31] ), .B(n95), .C(n94), .D(Packet_Out[31]), 
        .Z(n96) );
  OAI21M1P U244 ( .A(n373), .B(n12), .C(n96), .Z(n273) );
  OA21M1P U245 ( .A(n139), .B(n100), .C(Rst_n), .Z(n98) );
  ND2M1P U246 ( .A(n99), .B(n137), .Z(n138) );
  AOI21M1P U247 ( .A(n6), .B(n140), .C(n141), .Z(n132) );
  AOI22M1P U248 ( .A(\Queue[2][0] ), .B(n133), .C(\Queue[3][0] ), .D(n5), .Z(
        n101) );
  OAI21M1P U249 ( .A(n144), .B(n135), .C(n101), .Z(n272) );
  OAI21M1P U250 ( .A(n146), .B(n135), .C(n102), .Z(n271) );
  AOI22M1P U251 ( .A(\Queue[2][2] ), .B(n133), .C(n5), .D(\Queue[3][2] ), .Z(
        n103) );
  OAI21M1P U252 ( .A(n148), .B(n135), .C(n103), .Z(n270) );
  AOI22M1P U253 ( .A(\Queue[2][3] ), .B(n133), .C(n5), .D(\Queue[3][3] ), .Z(
        n104) );
  OAI21M1P U254 ( .A(n150), .B(n135), .C(n104), .Z(n269) );
  AOI22M1P U255 ( .A(\Queue[2][4] ), .B(n133), .C(n5), .D(\Queue[3][4] ), .Z(
        n105) );
  OAI21M1P U256 ( .A(n152), .B(n135), .C(n105), .Z(n268) );
  AOI22M1P U257 ( .A(\Queue[2][5] ), .B(n133), .C(n5), .D(\Queue[3][5] ), .Z(
        n106) );
  OAI21M1P U258 ( .A(n154), .B(n135), .C(n106), .Z(n267) );
  AOI22M1P U259 ( .A(\Queue[2][6] ), .B(n133), .C(n5), .D(\Queue[3][6] ), .Z(
        n107) );
  OAI21M1P U260 ( .A(n156), .B(n135), .C(n107), .Z(n266) );
  AOI22M1P U261 ( .A(\Queue[2][7] ), .B(n133), .C(n5), .D(\Queue[3][7] ), .Z(
        n108) );
  OAI21M1P U262 ( .A(n158), .B(n135), .C(n108), .Z(n265) );
  AOI22M1P U263 ( .A(\Queue[2][8] ), .B(n133), .C(n5), .D(\Queue[3][8] ), .Z(
        n109) );
  OAI21M1P U264 ( .A(n160), .B(n135), .C(n109), .Z(n264) );
  AOI22M1P U265 ( .A(\Queue[2][9] ), .B(n133), .C(n5), .D(\Queue[3][9] ), .Z(
        n110) );
  OAI21M1P U266 ( .A(n162), .B(n135), .C(n110), .Z(n263) );
  AOI22M1P U267 ( .A(\Queue[2][10] ), .B(n133), .C(n5), .D(\Queue[3][10] ), 
        .Z(n111) );
  OAI21M1P U268 ( .A(n164), .B(n135), .C(n111), .Z(n262) );
  AOI22M1P U269 ( .A(\Queue[2][11] ), .B(n133), .C(n5), .D(\Queue[3][11] ), 
        .Z(n112) );
  OAI21M1P U270 ( .A(n166), .B(n135), .C(n112), .Z(n261) );
  AOI22M1P U271 ( .A(\Queue[2][12] ), .B(n133), .C(n5), .D(\Queue[3][12] ), 
        .Z(n113) );
  OAI21M1P U272 ( .A(n168), .B(n135), .C(n113), .Z(n260) );
  AOI22M1P U273 ( .A(\Queue[2][13] ), .B(n133), .C(n5), .D(\Queue[3][13] ), 
        .Z(n114) );
  OAI21M1P U274 ( .A(n170), .B(n135), .C(n114), .Z(n259) );
  AOI22M1P U275 ( .A(\Queue[2][14] ), .B(n133), .C(n5), .D(\Queue[3][14] ), 
        .Z(n115) );
  OAI21M1P U276 ( .A(n172), .B(n135), .C(n115), .Z(n258) );
  AOI22M1P U277 ( .A(\Queue[2][15] ), .B(n133), .C(n5), .D(\Queue[3][15] ), 
        .Z(n116) );
  OAI21M1P U278 ( .A(n174), .B(n135), .C(n116), .Z(n257) );
  AOI22M1P U279 ( .A(\Queue[2][16] ), .B(n133), .C(n5), .D(\Queue[3][16] ), 
        .Z(n117) );
  OAI21M1P U280 ( .A(n176), .B(n135), .C(n117), .Z(n256) );
  AOI22M1P U281 ( .A(\Queue[2][17] ), .B(n133), .C(n5), .D(\Queue[3][17] ), 
        .Z(n118) );
  OAI21M1P U282 ( .A(n178), .B(n135), .C(n118), .Z(n255) );
  AOI22M1P U283 ( .A(\Queue[2][18] ), .B(n133), .C(n5), .D(\Queue[3][18] ), 
        .Z(n119) );
  OAI21M1P U284 ( .A(n180), .B(n135), .C(n119), .Z(n254) );
  AOI22M1P U285 ( .A(\Queue[2][19] ), .B(n133), .C(n5), .D(\Queue[3][19] ), 
        .Z(n120) );
  OAI21M1P U286 ( .A(n182), .B(n135), .C(n120), .Z(n253) );
  AOI22M1P U287 ( .A(\Queue[2][20] ), .B(n133), .C(n5), .D(\Queue[3][20] ), 
        .Z(n121) );
  OAI21M1P U288 ( .A(n184), .B(n135), .C(n121), .Z(n252) );
  AOI22M1P U289 ( .A(\Queue[2][21] ), .B(n133), .C(n5), .D(\Queue[3][21] ), 
        .Z(n122) );
  OAI21M1P U290 ( .A(n186), .B(n135), .C(n122), .Z(n251) );
  AOI22M1P U291 ( .A(\Queue[2][22] ), .B(n133), .C(n5), .D(\Queue[3][22] ), 
        .Z(n123) );
  OAI21M1P U292 ( .A(n188), .B(n135), .C(n123), .Z(n250) );
  AOI22M1P U293 ( .A(\Queue[2][23] ), .B(n133), .C(n5), .D(\Queue[3][23] ), 
        .Z(n124) );
  OAI21M1P U294 ( .A(n190), .B(n135), .C(n124), .Z(n249) );
  AOI22M1P U295 ( .A(\Queue[2][24] ), .B(n133), .C(n5), .D(\Queue[3][24] ), 
        .Z(n125) );
  OAI21M1P U296 ( .A(n192), .B(n135), .C(n125), .Z(n248) );
  AOI22M1P U297 ( .A(\Queue[2][25] ), .B(n133), .C(n5), .D(\Queue[3][25] ), 
        .Z(n126) );
  OAI21M1P U298 ( .A(n194), .B(n135), .C(n126), .Z(n247) );
  AOI22M1P U299 ( .A(\Queue[2][26] ), .B(n133), .C(n5), .D(\Queue[3][26] ), 
        .Z(n127) );
  OAI21M1P U300 ( .A(n196), .B(n135), .C(n127), .Z(n246) );
  AOI22M1P U301 ( .A(\Queue[2][27] ), .B(n133), .C(n5), .D(\Queue[3][27] ), 
        .Z(n128) );
  OAI21M1P U302 ( .A(n198), .B(n135), .C(n128), .Z(n245) );
  AOI22M1P U303 ( .A(\Queue[2][28] ), .B(n133), .C(n5), .D(\Queue[3][28] ), 
        .Z(n129) );
  OAI21M1P U304 ( .A(n200), .B(n135), .C(n129), .Z(n244) );
  AOI22M1P U305 ( .A(\Queue[2][29] ), .B(n133), .C(n5), .D(\Queue[3][29] ), 
        .Z(n130) );
  OAI21M1P U306 ( .A(n202), .B(n135), .C(n130), .Z(n243) );
  AOI22M1P U307 ( .A(\Queue[2][30] ), .B(n133), .C(n5), .D(\Queue[3][30] ), 
        .Z(n131) );
  OAI21M1P U308 ( .A(n204), .B(n135), .C(n131), .Z(n242) );
  AOI22M1P U309 ( .A(\Queue[2][31] ), .B(n133), .C(n5), .D(\Queue[3][31] ), 
        .Z(n134) );
  OAI21M1P U310 ( .A(n373), .B(n135), .C(n134), .Z(n241) );
  OA21M1P U311 ( .A(n139), .B(n140), .C(Rst_n), .Z(n136) );
  AOI21M1P U312 ( .A(n6), .B(n142), .C(n141), .Z(n205) );
  AOI22M1P U313 ( .A(\Queue[3][0] ), .B(n206), .C(n4), .D(\Queue[4][0] ), .Z(
        n143) );
  OAI21M1P U314 ( .A(n144), .B(n208), .C(n143), .Z(n240) );
  AOI22M1P U315 ( .A(\Queue[3][1] ), .B(n206), .C(n4), .D(\Queue[4][1] ), .Z(
        n145) );
  OAI21M1P U316 ( .A(n146), .B(n208), .C(n145), .Z(n239) );
  AOI22M1P U317 ( .A(\Queue[3][2] ), .B(n206), .C(n4), .D(\Queue[4][2] ), .Z(
        n147) );
  OAI21M1P U318 ( .A(n148), .B(n208), .C(n147), .Z(n238) );
  AOI22M1P U319 ( .A(\Queue[3][3] ), .B(n206), .C(n4), .D(\Queue[4][3] ), .Z(
        n149) );
  OAI21M1P U320 ( .A(n150), .B(n208), .C(n149), .Z(n237) );
  AOI22M1P U321 ( .A(\Queue[3][4] ), .B(n206), .C(n4), .D(\Queue[4][4] ), .Z(
        n151) );
  OAI21M1P U322 ( .A(n152), .B(n208), .C(n151), .Z(n236) );
  AOI22M1P U323 ( .A(\Queue[3][5] ), .B(n206), .C(n4), .D(\Queue[4][5] ), .Z(
        n153) );
  OAI21M1P U324 ( .A(n154), .B(n208), .C(n153), .Z(n235) );
  AOI22M1P U325 ( .A(\Queue[3][6] ), .B(n206), .C(n4), .D(\Queue[4][6] ), .Z(
        n155) );
  OAI21M1P U326 ( .A(n156), .B(n208), .C(n155), .Z(n234) );
  AOI22M1P U327 ( .A(\Queue[3][7] ), .B(n206), .C(n4), .D(\Queue[4][7] ), .Z(
        n157) );
  OAI21M1P U328 ( .A(n158), .B(n208), .C(n157), .Z(n233) );
  AOI22M1P U329 ( .A(\Queue[3][8] ), .B(n206), .C(n4), .D(\Queue[4][8] ), .Z(
        n159) );
  OAI21M1P U330 ( .A(n160), .B(n208), .C(n159), .Z(n232) );
  AOI22M1P U331 ( .A(\Queue[3][9] ), .B(n206), .C(n4), .D(\Queue[4][9] ), .Z(
        n161) );
  OAI21M1P U332 ( .A(n162), .B(n208), .C(n161), .Z(n231) );
  AOI22M1P U333 ( .A(\Queue[3][10] ), .B(n206), .C(n4), .D(\Queue[4][10] ), 
        .Z(n163) );
  OAI21M1P U334 ( .A(n164), .B(n208), .C(n163), .Z(n230) );
  AOI22M1P U335 ( .A(\Queue[3][11] ), .B(n206), .C(n4), .D(\Queue[4][11] ), 
        .Z(n165) );
  OAI21M1P U336 ( .A(n166), .B(n208), .C(n165), .Z(n229) );
  AOI22M1P U337 ( .A(\Queue[3][12] ), .B(n206), .C(n4), .D(\Queue[4][12] ), 
        .Z(n167) );
  OAI21M1P U338 ( .A(n168), .B(n208), .C(n167), .Z(n228) );
  AOI22M1P U339 ( .A(\Queue[3][13] ), .B(n206), .C(n4), .D(\Queue[4][13] ), 
        .Z(n169) );
  OAI21M1P U340 ( .A(n170), .B(n208), .C(n169), .Z(n227) );
  AOI22M1P U341 ( .A(\Queue[3][14] ), .B(n206), .C(n4), .D(\Queue[4][14] ), 
        .Z(n171) );
  OAI21M1P U342 ( .A(n172), .B(n208), .C(n171), .Z(n226) );
  AOI22M1P U343 ( .A(\Queue[3][15] ), .B(n206), .C(n4), .D(\Queue[4][15] ), 
        .Z(n173) );
  OAI21M1P U344 ( .A(n174), .B(n208), .C(n173), .Z(n225) );
  AOI22M1P U345 ( .A(\Queue[3][16] ), .B(n206), .C(n4), .D(\Queue[4][16] ), 
        .Z(n175) );
  OAI21M1P U346 ( .A(n176), .B(n208), .C(n175), .Z(n224) );
  AOI22M1P U347 ( .A(\Queue[3][17] ), .B(n206), .C(n4), .D(\Queue[4][17] ), 
        .Z(n177) );
  OAI21M1P U348 ( .A(n178), .B(n208), .C(n177), .Z(n223) );
  AOI22M1P U349 ( .A(\Queue[3][18] ), .B(n206), .C(n4), .D(\Queue[4][18] ), 
        .Z(n179) );
  OAI21M1P U350 ( .A(n180), .B(n208), .C(n179), .Z(n222) );
  AOI22M1P U351 ( .A(\Queue[3][19] ), .B(n206), .C(n4), .D(\Queue[4][19] ), 
        .Z(n181) );
  OAI21M1P U352 ( .A(n182), .B(n208), .C(n181), .Z(n221) );
  AOI22M1P U353 ( .A(\Queue[3][20] ), .B(n206), .C(n4), .D(\Queue[4][20] ), 
        .Z(n183) );
  OAI21M1P U354 ( .A(n184), .B(n208), .C(n183), .Z(n220) );
  AOI22M1P U355 ( .A(\Queue[3][21] ), .B(n206), .C(n4), .D(\Queue[4][21] ), 
        .Z(n185) );
  OAI21M1P U356 ( .A(n186), .B(n208), .C(n185), .Z(n219) );
  AOI22M1P U357 ( .A(\Queue[3][22] ), .B(n206), .C(n4), .D(\Queue[4][22] ), 
        .Z(n187) );
  OAI21M1P U358 ( .A(n188), .B(n208), .C(n187), .Z(n218) );
  AOI22M1P U359 ( .A(\Queue[3][23] ), .B(n206), .C(n4), .D(\Queue[4][23] ), 
        .Z(n189) );
  OAI21M1P U360 ( .A(n190), .B(n208), .C(n189), .Z(n217) );
  AOI22M1P U361 ( .A(\Queue[3][24] ), .B(n206), .C(n4), .D(\Queue[4][24] ), 
        .Z(n191) );
  OAI21M1P U362 ( .A(n192), .B(n208), .C(n191), .Z(n216) );
  AOI22M1P U363 ( .A(\Queue[3][25] ), .B(n206), .C(n4), .D(\Queue[4][25] ), 
        .Z(n193) );
  OAI21M1P U364 ( .A(n194), .B(n208), .C(n193), .Z(n215) );
  AOI22M1P U365 ( .A(\Queue[3][26] ), .B(n206), .C(n4), .D(\Queue[4][26] ), 
        .Z(n195) );
  OAI21M1P U366 ( .A(n196), .B(n208), .C(n195), .Z(n214) );
  AOI22M1P U367 ( .A(\Queue[3][27] ), .B(n206), .C(n4), .D(\Queue[4][27] ), 
        .Z(n197) );
  OAI21M1P U368 ( .A(n198), .B(n208), .C(n197), .Z(n213) );
  AOI22M1P U369 ( .A(\Queue[3][28] ), .B(n206), .C(n4), .D(\Queue[4][28] ), 
        .Z(n199) );
  OAI21M1P U370 ( .A(n200), .B(n208), .C(n199), .Z(n212) );
  AOI22M1P U371 ( .A(\Queue[3][29] ), .B(n206), .C(n4), .D(\Queue[4][29] ), 
        .Z(n201) );
  OAI21M1P U372 ( .A(n202), .B(n208), .C(n201), .Z(n211) );
  AOI22M1P U373 ( .A(\Queue[3][30] ), .B(n206), .C(n4), .D(\Queue[4][30] ), 
        .Z(n203) );
  OAI21M1P U374 ( .A(n204), .B(n208), .C(n203), .Z(n210) );
  AOI22M1P U375 ( .A(\Queue[3][31] ), .B(n206), .C(n4), .D(\Queue[4][31] ), 
        .Z(n207) );
  OAI21M1P U376 ( .A(n373), .B(n208), .C(n207), .Z(n209) );
  N1M1P U377 ( .A(n2), .Z(Empty) );
  AOI22M1P U378 ( .A(n376), .B(n375), .C(n374), .D(Empty), .Z(n1) );
endmodule


module Packet_Queue_9 ( Clk_r, Rst_n, Packet_In, Read_Ack, Write_Ack, 
        Packet_Out, Empty, Full );
  input [31:0] Packet_In;
  output [31:0] Packet_Out;
  input Clk_r, Rst_n, Read_Ack, Write_Ack;
  output Empty, Full;
  wire   \Queue[4][31] , \Queue[4][30] , \Queue[4][29] , \Queue[4][28] ,
         \Queue[4][27] , \Queue[4][26] , \Queue[4][25] , \Queue[4][24] ,
         \Queue[4][23] , \Queue[4][22] , \Queue[4][21] , \Queue[4][20] ,
         \Queue[4][19] , \Queue[4][18] , \Queue[4][17] , \Queue[4][16] ,
         \Queue[4][15] , \Queue[4][14] , \Queue[4][13] , \Queue[4][12] ,
         \Queue[4][11] , \Queue[4][10] , \Queue[4][9] , \Queue[4][8] ,
         \Queue[4][7] , \Queue[4][6] , \Queue[4][5] , \Queue[4][4] ,
         \Queue[4][3] , \Queue[4][2] , \Queue[4][1] , \Queue[4][0] ,
         \Queue[3][31] , \Queue[3][30] , \Queue[3][29] , \Queue[3][28] ,
         \Queue[3][27] , \Queue[3][26] , \Queue[3][25] , \Queue[3][24] ,
         \Queue[3][23] , \Queue[3][22] , \Queue[3][21] , \Queue[3][20] ,
         \Queue[3][19] , \Queue[3][18] , \Queue[3][17] , \Queue[3][16] ,
         \Queue[3][15] , \Queue[3][14] , \Queue[3][13] , \Queue[3][12] ,
         \Queue[3][11] , \Queue[3][10] , \Queue[3][9] , \Queue[3][8] ,
         \Queue[3][7] , \Queue[3][6] , \Queue[3][5] , \Queue[3][4] ,
         \Queue[3][3] , \Queue[3][2] , \Queue[3][1] , \Queue[3][0] ,
         \Queue[2][31] , \Queue[2][30] , \Queue[2][29] , \Queue[2][28] ,
         \Queue[2][27] , \Queue[2][26] , \Queue[2][25] , \Queue[2][24] ,
         \Queue[2][23] , \Queue[2][22] , \Queue[2][21] , \Queue[2][20] ,
         \Queue[2][19] , \Queue[2][18] , \Queue[2][17] , \Queue[2][16] ,
         \Queue[2][15] , \Queue[2][14] , \Queue[2][13] , \Queue[2][12] ,
         \Queue[2][11] , \Queue[2][10] , \Queue[2][9] , \Queue[2][8] ,
         \Queue[2][7] , \Queue[2][6] , \Queue[2][5] , \Queue[2][4] ,
         \Queue[2][3] , \Queue[2][2] , \Queue[2][1] , \Queue[2][0] ,
         \Queue[1][31] , \Queue[1][30] , \Queue[1][29] , \Queue[1][28] ,
         \Queue[1][27] , \Queue[1][26] , \Queue[1][25] , \Queue[1][24] ,
         \Queue[1][23] , \Queue[1][22] , \Queue[1][21] , \Queue[1][20] ,
         \Queue[1][19] , \Queue[1][18] , \Queue[1][17] , \Queue[1][16] ,
         \Queue[1][15] , \Queue[1][14] , \Queue[1][13] , \Queue[1][12] ,
         \Queue[1][11] , \Queue[1][10] , \Queue[1][9] , \Queue[1][8] ,
         \Queue[1][7] , \Queue[1][6] , \Queue[1][5] , \Queue[1][4] ,
         \Queue[1][3] , \Queue[1][2] , \Queue[1][1] , \Queue[1][0] , n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546;
  wire   [2:0] Count;

  FDN2QM1P \Count_reg[0]  ( .D(n381), .CPN(Clk_r), .CD(Rst_n), .Q(Count[0]) );
  FDN2QM1P \Count_reg[1]  ( .D(n382), .CPN(Clk_r), .CD(Rst_n), .Q(Count[1]) );
  FDN2QM1P \Count_reg[2]  ( .D(n383), .CPN(Clk_r), .CD(Rst_n), .Q(Count[2]) );
  FDN1QM1P \Queue_reg[4][30]  ( .D(n415), .CPN(Clk_r), .Q(\Queue[4][30] ) );
  FDN1QM1P \Queue_reg[3][30]  ( .D(n543), .CPN(Clk_r), .Q(\Queue[3][30] ) );
  FDN1QM1P \Queue_reg[2][30]  ( .D(n511), .CPN(Clk_r), .Q(\Queue[2][30] ) );
  FDN1QM1P \Queue_reg[4][29]  ( .D(n414), .CPN(Clk_r), .Q(\Queue[4][29] ) );
  FDN1QM1P \Queue_reg[3][29]  ( .D(n542), .CPN(Clk_r), .Q(\Queue[3][29] ) );
  FDN1QM1P \Queue_reg[2][29]  ( .D(n510), .CPN(Clk_r), .Q(\Queue[2][29] ) );
  FDN1QM1P \Queue_reg[4][28]  ( .D(n413), .CPN(Clk_r), .Q(\Queue[4][28] ) );
  FDN1QM1P \Queue_reg[3][28]  ( .D(n541), .CPN(Clk_r), .Q(\Queue[3][28] ) );
  FDN1QM1P \Queue_reg[2][28]  ( .D(n509), .CPN(Clk_r), .Q(\Queue[2][28] ) );
  FDN1QM1P \Queue_reg[4][27]  ( .D(n412), .CPN(Clk_r), .Q(\Queue[4][27] ) );
  FDN1QM1P \Queue_reg[3][27]  ( .D(n540), .CPN(Clk_r), .Q(\Queue[3][27] ) );
  FDN1QM1P \Queue_reg[2][27]  ( .D(n508), .CPN(Clk_r), .Q(\Queue[2][27] ) );
  FDN1QM1P \Queue_reg[4][26]  ( .D(n411), .CPN(Clk_r), .Q(\Queue[4][26] ) );
  FDN1QM1P \Queue_reg[3][26]  ( .D(n539), .CPN(Clk_r), .Q(\Queue[3][26] ) );
  FDN1QM1P \Queue_reg[2][26]  ( .D(n507), .CPN(Clk_r), .Q(\Queue[2][26] ) );
  FDN1QM1P \Queue_reg[4][25]  ( .D(n410), .CPN(Clk_r), .Q(\Queue[4][25] ) );
  FDN1QM1P \Queue_reg[3][25]  ( .D(n538), .CPN(Clk_r), .Q(\Queue[3][25] ) );
  FDN1QM1P \Queue_reg[2][25]  ( .D(n506), .CPN(Clk_r), .Q(\Queue[2][25] ) );
  FDN1QM1P \Queue_reg[4][24]  ( .D(n409), .CPN(Clk_r), .Q(\Queue[4][24] ) );
  FDN1QM1P \Queue_reg[3][24]  ( .D(n537), .CPN(Clk_r), .Q(\Queue[3][24] ) );
  FDN1QM1P \Queue_reg[2][24]  ( .D(n505), .CPN(Clk_r), .Q(\Queue[2][24] ) );
  FDN1QM1P \Queue_reg[4][23]  ( .D(n408), .CPN(Clk_r), .Q(\Queue[4][23] ) );
  FDN1QM1P \Queue_reg[3][23]  ( .D(n536), .CPN(Clk_r), .Q(\Queue[3][23] ) );
  FDN1QM1P \Queue_reg[2][23]  ( .D(n504), .CPN(Clk_r), .Q(\Queue[2][23] ) );
  FDN1QM1P \Queue_reg[4][22]  ( .D(n407), .CPN(Clk_r), .Q(\Queue[4][22] ) );
  FDN1QM1P \Queue_reg[3][22]  ( .D(n535), .CPN(Clk_r), .Q(\Queue[3][22] ) );
  FDN1QM1P \Queue_reg[2][22]  ( .D(n503), .CPN(Clk_r), .Q(\Queue[2][22] ) );
  FDN1QM1P \Queue_reg[4][21]  ( .D(n406), .CPN(Clk_r), .Q(\Queue[4][21] ) );
  FDN1QM1P \Queue_reg[3][21]  ( .D(n534), .CPN(Clk_r), .Q(\Queue[3][21] ) );
  FDN1QM1P \Queue_reg[2][21]  ( .D(n502), .CPN(Clk_r), .Q(\Queue[2][21] ) );
  FDN1QM1P \Queue_reg[4][20]  ( .D(n405), .CPN(Clk_r), .Q(\Queue[4][20] ) );
  FDN1QM1P \Queue_reg[3][20]  ( .D(n533), .CPN(Clk_r), .Q(\Queue[3][20] ) );
  FDN1QM1P \Queue_reg[2][20]  ( .D(n501), .CPN(Clk_r), .Q(\Queue[2][20] ) );
  FDN1QM1P \Queue_reg[4][19]  ( .D(n404), .CPN(Clk_r), .Q(\Queue[4][19] ) );
  FDN1QM1P \Queue_reg[3][19]  ( .D(n532), .CPN(Clk_r), .Q(\Queue[3][19] ) );
  FDN1QM1P \Queue_reg[2][19]  ( .D(n500), .CPN(Clk_r), .Q(\Queue[2][19] ) );
  FDN1QM1P \Queue_reg[4][18]  ( .D(n403), .CPN(Clk_r), .Q(\Queue[4][18] ) );
  FDN1QM1P \Queue_reg[3][18]  ( .D(n531), .CPN(Clk_r), .Q(\Queue[3][18] ) );
  FDN1QM1P \Queue_reg[2][18]  ( .D(n499), .CPN(Clk_r), .Q(\Queue[2][18] ) );
  FDN1QM1P \Queue_reg[4][17]  ( .D(n402), .CPN(Clk_r), .Q(\Queue[4][17] ) );
  FDN1QM1P \Queue_reg[3][17]  ( .D(n530), .CPN(Clk_r), .Q(\Queue[3][17] ) );
  FDN1QM1P \Queue_reg[2][17]  ( .D(n498), .CPN(Clk_r), .Q(\Queue[2][17] ) );
  FDN1QM1P \Queue_reg[4][16]  ( .D(n401), .CPN(Clk_r), .Q(\Queue[4][16] ) );
  FDN1QM1P \Queue_reg[3][16]  ( .D(n529), .CPN(Clk_r), .Q(\Queue[3][16] ) );
  FDN1QM1P \Queue_reg[2][16]  ( .D(n497), .CPN(Clk_r), .Q(\Queue[2][16] ) );
  FDN1QM1P \Queue_reg[4][15]  ( .D(n400), .CPN(Clk_r), .Q(\Queue[4][15] ) );
  FDN1QM1P \Queue_reg[3][15]  ( .D(n528), .CPN(Clk_r), .Q(\Queue[3][15] ) );
  FDN1QM1P \Queue_reg[2][15]  ( .D(n496), .CPN(Clk_r), .Q(\Queue[2][15] ) );
  FDN1QM1P \Queue_reg[4][14]  ( .D(n399), .CPN(Clk_r), .Q(\Queue[4][14] ) );
  FDN1QM1P \Queue_reg[3][14]  ( .D(n527), .CPN(Clk_r), .Q(\Queue[3][14] ) );
  FDN1QM1P \Queue_reg[2][14]  ( .D(n495), .CPN(Clk_r), .Q(\Queue[2][14] ) );
  FDN1QM1P \Queue_reg[4][13]  ( .D(n398), .CPN(Clk_r), .Q(\Queue[4][13] ) );
  FDN1QM1P \Queue_reg[3][13]  ( .D(n526), .CPN(Clk_r), .Q(\Queue[3][13] ) );
  FDN1QM1P \Queue_reg[2][13]  ( .D(n494), .CPN(Clk_r), .Q(\Queue[2][13] ) );
  FDN1QM1P \Queue_reg[4][12]  ( .D(n397), .CPN(Clk_r), .Q(\Queue[4][12] ) );
  FDN1QM1P \Queue_reg[3][12]  ( .D(n525), .CPN(Clk_r), .Q(\Queue[3][12] ) );
  FDN1QM1P \Queue_reg[2][12]  ( .D(n493), .CPN(Clk_r), .Q(\Queue[2][12] ) );
  FDN1QM1P \Queue_reg[4][11]  ( .D(n396), .CPN(Clk_r), .Q(\Queue[4][11] ) );
  FDN1QM1P \Queue_reg[3][11]  ( .D(n524), .CPN(Clk_r), .Q(\Queue[3][11] ) );
  FDN1QM1P \Queue_reg[2][11]  ( .D(n492), .CPN(Clk_r), .Q(\Queue[2][11] ) );
  FDN1QM1P \Queue_reg[4][10]  ( .D(n395), .CPN(Clk_r), .Q(\Queue[4][10] ) );
  FDN1QM1P \Queue_reg[3][10]  ( .D(n523), .CPN(Clk_r), .Q(\Queue[3][10] ) );
  FDN1QM1P \Queue_reg[2][10]  ( .D(n491), .CPN(Clk_r), .Q(\Queue[2][10] ) );
  FDN1QM1P \Queue_reg[4][9]  ( .D(n394), .CPN(Clk_r), .Q(\Queue[4][9] ) );
  FDN1QM1P \Queue_reg[3][9]  ( .D(n522), .CPN(Clk_r), .Q(\Queue[3][9] ) );
  FDN1QM1P \Queue_reg[2][9]  ( .D(n490), .CPN(Clk_r), .Q(\Queue[2][9] ) );
  FDN1QM1P \Queue_reg[4][8]  ( .D(n393), .CPN(Clk_r), .Q(\Queue[4][8] ) );
  FDN1QM1P \Queue_reg[3][8]  ( .D(n521), .CPN(Clk_r), .Q(\Queue[3][8] ) );
  FDN1QM1P \Queue_reg[2][8]  ( .D(n489), .CPN(Clk_r), .Q(\Queue[2][8] ) );
  FDN1QM1P \Queue_reg[4][7]  ( .D(n392), .CPN(Clk_r), .Q(\Queue[4][7] ) );
  FDN1QM1P \Queue_reg[3][7]  ( .D(n520), .CPN(Clk_r), .Q(\Queue[3][7] ) );
  FDN1QM1P \Queue_reg[2][7]  ( .D(n488), .CPN(Clk_r), .Q(\Queue[2][7] ) );
  FDN1QM1P \Queue_reg[4][6]  ( .D(n391), .CPN(Clk_r), .Q(\Queue[4][6] ) );
  FDN1QM1P \Queue_reg[3][6]  ( .D(n519), .CPN(Clk_r), .Q(\Queue[3][6] ) );
  FDN1QM1P \Queue_reg[2][6]  ( .D(n487), .CPN(Clk_r), .Q(\Queue[2][6] ) );
  FDN1QM1P \Queue_reg[4][5]  ( .D(n390), .CPN(Clk_r), .Q(\Queue[4][5] ) );
  FDN1QM1P \Queue_reg[3][5]  ( .D(n518), .CPN(Clk_r), .Q(\Queue[3][5] ) );
  FDN1QM1P \Queue_reg[2][5]  ( .D(n486), .CPN(Clk_r), .Q(\Queue[2][5] ) );
  FDN1QM1P \Queue_reg[4][4]  ( .D(n389), .CPN(Clk_r), .Q(\Queue[4][4] ) );
  FDN1QM1P \Queue_reg[3][4]  ( .D(n517), .CPN(Clk_r), .Q(\Queue[3][4] ) );
  FDN1QM1P \Queue_reg[2][4]  ( .D(n485), .CPN(Clk_r), .Q(\Queue[2][4] ) );
  FDN1QM1P \Queue_reg[4][3]  ( .D(n388), .CPN(Clk_r), .Q(\Queue[4][3] ) );
  FDN1QM1P \Queue_reg[3][3]  ( .D(n516), .CPN(Clk_r), .Q(\Queue[3][3] ) );
  FDN1QM1P \Queue_reg[2][3]  ( .D(n484), .CPN(Clk_r), .Q(\Queue[2][3] ) );
  FDN1QM1P \Queue_reg[4][2]  ( .D(n387), .CPN(Clk_r), .Q(\Queue[4][2] ) );
  FDN1QM1P \Queue_reg[3][2]  ( .D(n515), .CPN(Clk_r), .Q(\Queue[3][2] ) );
  FDN1QM1P \Queue_reg[2][2]  ( .D(n483), .CPN(Clk_r), .Q(\Queue[2][2] ) );
  FDN1QM1P \Queue_reg[4][1]  ( .D(n386), .CPN(Clk_r), .Q(\Queue[4][1] ) );
  FDN1QM1P \Queue_reg[3][1]  ( .D(n514), .CPN(Clk_r), .Q(\Queue[3][1] ) );
  FDN1QM1P \Queue_reg[2][1]  ( .D(n482), .CPN(Clk_r), .Q(\Queue[2][1] ) );
  FDN1QM1P \Queue_reg[4][0]  ( .D(n385), .CPN(Clk_r), .Q(\Queue[4][0] ) );
  FDN1QM1P \Queue_reg[3][0]  ( .D(n513), .CPN(Clk_r), .Q(\Queue[3][0] ) );
  FDN1QM1P \Queue_reg[2][0]  ( .D(n481), .CPN(Clk_r), .Q(\Queue[2][0] ) );
  FDN1QM1P \Queue_reg[4][31]  ( .D(n384), .CPN(Clk_r), .Q(\Queue[4][31] ) );
  FDN1QM1P \Queue_reg[3][31]  ( .D(n544), .CPN(Clk_r), .Q(\Queue[3][31] ) );
  FDN1QM1P \Queue_reg[2][31]  ( .D(n512), .CPN(Clk_r), .Q(\Queue[2][31] ) );
  FDN2QM1P Full_reg ( .D(n416), .CPN(Clk_r), .CD(Rst_n), .Q(Full) );
  FDN1QM1P \Queue_reg[1][31]  ( .D(n448), .CPN(Clk_r), .Q(\Queue[1][31] ) );
  FDN1QM1P \Queue_reg[0][31]  ( .D(n480), .CPN(Clk_r), .Q(Packet_Out[31]) );
  FDN1QM1P \Queue_reg[1][30]  ( .D(n447), .CPN(Clk_r), .Q(\Queue[1][30] ) );
  FDN1QM1P \Queue_reg[0][30]  ( .D(n479), .CPN(Clk_r), .Q(Packet_Out[30]) );
  FDN1QM1P \Queue_reg[1][29]  ( .D(n446), .CPN(Clk_r), .Q(\Queue[1][29] ) );
  FDN1QM1P \Queue_reg[0][29]  ( .D(n478), .CPN(Clk_r), .Q(Packet_Out[29]) );
  FDN1QM1P \Queue_reg[1][28]  ( .D(n445), .CPN(Clk_r), .Q(\Queue[1][28] ) );
  FDN1QM1P \Queue_reg[0][28]  ( .D(n477), .CPN(Clk_r), .Q(Packet_Out[28]) );
  FDN1QM1P \Queue_reg[1][27]  ( .D(n444), .CPN(Clk_r), .Q(\Queue[1][27] ) );
  FDN1QM1P \Queue_reg[0][27]  ( .D(n476), .CPN(Clk_r), .Q(Packet_Out[27]) );
  FDN1QM1P \Queue_reg[1][26]  ( .D(n443), .CPN(Clk_r), .Q(\Queue[1][26] ) );
  FDN1QM1P \Queue_reg[0][26]  ( .D(n475), .CPN(Clk_r), .Q(Packet_Out[26]) );
  FDN1QM1P \Queue_reg[1][25]  ( .D(n442), .CPN(Clk_r), .Q(\Queue[1][25] ) );
  FDN1QM1P \Queue_reg[0][25]  ( .D(n474), .CPN(Clk_r), .Q(Packet_Out[25]) );
  FDN1QM1P \Queue_reg[1][24]  ( .D(n441), .CPN(Clk_r), .Q(\Queue[1][24] ) );
  FDN1QM1P \Queue_reg[0][24]  ( .D(n473), .CPN(Clk_r), .Q(Packet_Out[24]) );
  FDN1QM1P \Queue_reg[1][23]  ( .D(n440), .CPN(Clk_r), .Q(\Queue[1][23] ) );
  FDN1QM1P \Queue_reg[0][23]  ( .D(n472), .CPN(Clk_r), .Q(Packet_Out[23]) );
  FDN1QM1P \Queue_reg[1][22]  ( .D(n439), .CPN(Clk_r), .Q(\Queue[1][22] ) );
  FDN1QM1P \Queue_reg[0][22]  ( .D(n471), .CPN(Clk_r), .Q(Packet_Out[22]) );
  FDN1QM1P \Queue_reg[1][21]  ( .D(n438), .CPN(Clk_r), .Q(\Queue[1][21] ) );
  FDN1QM1P \Queue_reg[0][21]  ( .D(n470), .CPN(Clk_r), .Q(Packet_Out[21]) );
  FDN1QM1P \Queue_reg[1][20]  ( .D(n437), .CPN(Clk_r), .Q(\Queue[1][20] ) );
  FDN1QM1P \Queue_reg[0][20]  ( .D(n469), .CPN(Clk_r), .Q(Packet_Out[20]) );
  FDN1QM1P \Queue_reg[1][19]  ( .D(n436), .CPN(Clk_r), .Q(\Queue[1][19] ) );
  FDN1QM1P \Queue_reg[0][19]  ( .D(n468), .CPN(Clk_r), .Q(Packet_Out[19]) );
  FDN1QM1P \Queue_reg[1][18]  ( .D(n435), .CPN(Clk_r), .Q(\Queue[1][18] ) );
  FDN1QM1P \Queue_reg[0][18]  ( .D(n467), .CPN(Clk_r), .Q(Packet_Out[18]) );
  FDN1QM1P \Queue_reg[1][17]  ( .D(n434), .CPN(Clk_r), .Q(\Queue[1][17] ) );
  FDN1QM1P \Queue_reg[0][17]  ( .D(n466), .CPN(Clk_r), .Q(Packet_Out[17]) );
  FDN1QM1P \Queue_reg[1][16]  ( .D(n433), .CPN(Clk_r), .Q(\Queue[1][16] ) );
  FDN1QM1P \Queue_reg[0][16]  ( .D(n465), .CPN(Clk_r), .Q(Packet_Out[16]) );
  FDN1QM1P \Queue_reg[1][15]  ( .D(n432), .CPN(Clk_r), .Q(\Queue[1][15] ) );
  FDN1QM1P \Queue_reg[0][15]  ( .D(n464), .CPN(Clk_r), .Q(Packet_Out[15]) );
  FDN1QM1P \Queue_reg[1][14]  ( .D(n431), .CPN(Clk_r), .Q(\Queue[1][14] ) );
  FDN1QM1P \Queue_reg[0][14]  ( .D(n463), .CPN(Clk_r), .Q(Packet_Out[14]) );
  FDN1QM1P \Queue_reg[1][13]  ( .D(n430), .CPN(Clk_r), .Q(\Queue[1][13] ) );
  FDN1QM1P \Queue_reg[0][13]  ( .D(n462), .CPN(Clk_r), .Q(Packet_Out[13]) );
  FDN1QM1P \Queue_reg[1][12]  ( .D(n429), .CPN(Clk_r), .Q(\Queue[1][12] ) );
  FDN1QM1P \Queue_reg[0][12]  ( .D(n461), .CPN(Clk_r), .Q(Packet_Out[12]) );
  FDN1QM1P \Queue_reg[1][11]  ( .D(n428), .CPN(Clk_r), .Q(\Queue[1][11] ) );
  FDN1QM1P \Queue_reg[0][11]  ( .D(n460), .CPN(Clk_r), .Q(Packet_Out[11]) );
  FDN1QM1P \Queue_reg[1][10]  ( .D(n427), .CPN(Clk_r), .Q(\Queue[1][10] ) );
  FDN1QM1P \Queue_reg[0][10]  ( .D(n459), .CPN(Clk_r), .Q(Packet_Out[10]) );
  FDN1QM1P \Queue_reg[1][9]  ( .D(n426), .CPN(Clk_r), .Q(\Queue[1][9] ) );
  FDN1QM1P \Queue_reg[0][9]  ( .D(n458), .CPN(Clk_r), .Q(Packet_Out[9]) );
  FDN1QM1P \Queue_reg[1][8]  ( .D(n425), .CPN(Clk_r), .Q(\Queue[1][8] ) );
  FDN1QM1P \Queue_reg[0][8]  ( .D(n457), .CPN(Clk_r), .Q(Packet_Out[8]) );
  FDN1QM1P \Queue_reg[1][7]  ( .D(n424), .CPN(Clk_r), .Q(\Queue[1][7] ) );
  FDN1QM1P \Queue_reg[0][7]  ( .D(n456), .CPN(Clk_r), .Q(Packet_Out[7]) );
  FDN1QM1P \Queue_reg[1][6]  ( .D(n423), .CPN(Clk_r), .Q(\Queue[1][6] ) );
  FDN1QM1P \Queue_reg[0][6]  ( .D(n455), .CPN(Clk_r), .Q(Packet_Out[6]) );
  FDN1QM1P \Queue_reg[1][5]  ( .D(n422), .CPN(Clk_r), .Q(\Queue[1][5] ) );
  FDN1QM1P \Queue_reg[0][5]  ( .D(n454), .CPN(Clk_r), .Q(Packet_Out[5]) );
  FDN1QM1P \Queue_reg[1][4]  ( .D(n421), .CPN(Clk_r), .Q(\Queue[1][4] ) );
  FDN1QM1P \Queue_reg[0][4]  ( .D(n453), .CPN(Clk_r), .Q(Packet_Out[4]) );
  FDN1QM1P \Queue_reg[1][3]  ( .D(n420), .CPN(Clk_r), .Q(\Queue[1][3] ) );
  FDN1QM1P \Queue_reg[0][3]  ( .D(n452), .CPN(Clk_r), .Q(Packet_Out[3]) );
  FDN1QM1P \Queue_reg[1][2]  ( .D(n419), .CPN(Clk_r), .Q(\Queue[1][2] ) );
  FDN1QM1P \Queue_reg[0][2]  ( .D(n451), .CPN(Clk_r), .Q(Packet_Out[2]) );
  FDN1QM1P \Queue_reg[1][1]  ( .D(n418), .CPN(Clk_r), .Q(\Queue[1][1] ) );
  FDN1QM1P \Queue_reg[0][1]  ( .D(n450), .CPN(Clk_r), .Q(Packet_Out[1]) );
  FDN1QM1P \Queue_reg[1][0]  ( .D(n417), .CPN(Clk_r), .Q(\Queue[1][0] ) );
  FDN1QM1P \Queue_reg[0][0]  ( .D(n449), .CPN(Clk_r), .Q(Packet_Out[0]) );
  FDN2QM1P Empty_reg ( .D(n546), .CPN(Clk_r), .CD(Rst_n), .Q(n545) );
  NR3M1P U3 ( .A(Count[0]), .B(Count[2]), .C(n26), .Z(n104) );
  BUFM1P U4 ( .A(n63), .Z(n9) );
  BUFM1P U5 ( .A(n101), .Z(n11) );
  N1M2P U6 ( .A(n66), .Z(n98) );
  BUFM2P U7 ( .A(n63), .Z(n8) );
  BUFM1P U8 ( .A(n136), .Z(n12) );
  BUFM1P U9 ( .A(n137), .Z(n14) );
  BUFM1P U10 ( .A(n374), .Z(n16) );
  BUFM2P U11 ( .A(n137), .Z(n13) );
  BUFM2P U12 ( .A(n136), .Z(n3) );
  BUFM2P U13 ( .A(n374), .Z(n15) );
  N1M1P U14 ( .A(Read_Ack), .Z(n141) );
  ND2M1P U15 ( .A(Read_Ack), .B(Rst_n), .Z(n145) );
  NR3M1P U16 ( .A(Count[2]), .B(n27), .C(n26), .Z(n144) );
  NR3M1P U17 ( .A(n27), .B(Count[2]), .C(Count[1]), .Z(n380) );
  OAI211M4P U18 ( .A(n144), .B(n141), .C(Write_Ack), .D(n102), .Z(n139) );
  NR2FM3P U19 ( .A(n65), .B(n25), .Z(n24) );
  AOI21M3P U20 ( .A(Write_Ack), .B(n380), .C(n145), .Z(n99) );
  OAI211M4P U21 ( .A(n146), .B(n141), .C(Write_Ack), .D(n140), .Z(n376) );
  OAI21M2P U22 ( .A(Write_Ack), .B(Read_Ack), .C(n28), .Z(n60) );
  NR2M3P U23 ( .A(Read_Ack), .B(n103), .Z(n22) );
  NR3M1P U24 ( .A(Count[0]), .B(Count[1]), .C(n23), .Z(n146) );
  N1M1P U25 ( .A(Count[0]), .Z(n27) );
  N1M1P U26 ( .A(Count[1]), .Z(n26) );
  N1M1P U27 ( .A(Count[2]), .Z(n23) );
  OAI21M1P U28 ( .A(n65), .B(n64), .C(n145), .Z(n66) );
  AOI21M6P U29 ( .A(Write_Ack), .B(n104), .C(n145), .Z(n61) );
  ND2M2P U30 ( .A(n22), .B(Rst_n), .Z(n65) );
  N1M1P U31 ( .A(Packet_In[27]), .Z(n202) );
  N1M1P U32 ( .A(Packet_In[28]), .Z(n204) );
  N1M1P U33 ( .A(Packet_In[30]), .Z(n208) );
  N1M1P U34 ( .A(Packet_In[23]), .Z(n194) );
  N1M1P U35 ( .A(Packet_In[25]), .Z(n198) );
  N1M1P U36 ( .A(Packet_In[26]), .Z(n200) );
  N1M1P U37 ( .A(Packet_In[29]), .Z(n206) );
  N1M1P U38 ( .A(Packet_In[31]), .Z(n377) );
  N1M1P U39 ( .A(Packet_In[0]), .Z(n148) );
  N1M1P U40 ( .A(Packet_In[24]), .Z(n196) );
  N1M1P U41 ( .A(Packet_In[22]), .Z(n192) );
  N1M1P U42 ( .A(Packet_In[6]), .Z(n160) );
  N1M1P U43 ( .A(Packet_In[2]), .Z(n152) );
  N1M1P U44 ( .A(Packet_In[4]), .Z(n156) );
  N1M1P U45 ( .A(Packet_In[8]), .Z(n164) );
  N1M1P U46 ( .A(Packet_In[5]), .Z(n158) );
  N1M1P U47 ( .A(Packet_In[3]), .Z(n154) );
  N1M1P U48 ( .A(Packet_In[9]), .Z(n166) );
  N1M1P U49 ( .A(Packet_In[7]), .Z(n162) );
  N1M1P U50 ( .A(Packet_In[1]), .Z(n150) );
  N1M1P U51 ( .A(Packet_In[10]), .Z(n168) );
  N1M1P U52 ( .A(Packet_In[11]), .Z(n170) );
  N1M1P U53 ( .A(Packet_In[19]), .Z(n186) );
  N1M1P U54 ( .A(Packet_In[18]), .Z(n184) );
  N1M1P U55 ( .A(Packet_In[13]), .Z(n174) );
  N1M1P U56 ( .A(Packet_In[20]), .Z(n188) );
  N1M1P U57 ( .A(Packet_In[12]), .Z(n172) );
  N1M1P U58 ( .A(Packet_In[17]), .Z(n182) );
  N1M1P U59 ( .A(Packet_In[21]), .Z(n190) );
  N1M1P U60 ( .A(Packet_In[15]), .Z(n178) );
  N1M1P U61 ( .A(Packet_In[16]), .Z(n180) );
  N1M1P U62 ( .A(Packet_In[14]), .Z(n176) );
  BUFM4P U63 ( .A(n101), .Z(n10) );
  OAI211M1P U64 ( .A(n380), .B(n141), .C(Write_Ack), .D(n66), .Z(n101) );
  BUFM2P U65 ( .A(n61), .Z(n6) );
  AOI21M6P U66 ( .A(Write_Ack), .B(n146), .C(n145), .Z(n373) );
  BUFM2P U67 ( .A(n60), .Z(n5) );
  BUFM2P U68 ( .A(n60), .Z(n4) );
  BUFM2P U69 ( .A(n61), .Z(n7) );
  OAI211M1P U70 ( .A(n104), .B(n141), .C(Write_Ack), .D(n28), .Z(n63) );
  N1M2P U71 ( .A(n22), .Z(n143) );
  N1M2P U72 ( .A(Write_Ack), .Z(n103) );
  AOI22CDNM1P U73 ( .A(n21), .B(n27), .C(n27), .D(n22), .Z(n18) );
  OA21M1P U74 ( .A(n143), .B(n144), .C(Rst_n), .Z(n140) );
  OA21M1P U75 ( .A(n143), .B(n380), .C(Rst_n), .Z(n28) );
  OA21M1P U76 ( .A(n143), .B(n104), .C(Rst_n), .Z(n102) );
  OAI211M1P U77 ( .A(n104), .B(n143), .C(Rst_n), .D(n142), .Z(n137) );
  OAI211M1P U78 ( .A(n144), .B(n143), .C(Rst_n), .D(n142), .Z(n374) );
  NR2M1P U79 ( .A(n141), .B(Write_Ack), .Z(n379) );
  NR2M1P U80 ( .A(n22), .B(n379), .Z(n378) );
  AOI22CDNM1P U81 ( .A(n378), .B(n27), .C(n378), .D(n27), .Z(n381) );
  N1M1P U82 ( .A(n379), .Z(n21) );
  AOI22CDNM1P U83 ( .A(Count[1]), .B(n18), .C(n18), .D(Count[1]), .Z(n382) );
  ND3M1P U84 ( .A(n27), .B(n23), .C(n26), .Z(n64) );
  ND2M1P U85 ( .A(Count[1]), .B(Read_Ack), .Z(n17) );
  OAI211M1P U86 ( .A(Count[1]), .B(n143), .C(n18), .D(n17), .Z(n19) );
  AOI22M1P U87 ( .A(n22), .B(n144), .C(Count[2]), .D(n19), .Z(n20) );
  OAI21M1P U88 ( .A(n64), .B(n21), .C(n20), .Z(n383) );
  N1M1P U89 ( .A(n146), .Z(n25) );
  AOI22CDNM1P U90 ( .A(n24), .B(n377), .C(\Queue[4][31] ), .D(n24), .Z(n384)
         );
  AOI22CDNM1P U91 ( .A(n24), .B(n148), .C(\Queue[4][0] ), .D(n24), .Z(n385) );
  AOI22CDNM1P U92 ( .A(n24), .B(n150), .C(\Queue[4][1] ), .D(n24), .Z(n386) );
  AOI22CDNM1P U93 ( .A(n24), .B(n152), .C(\Queue[4][2] ), .D(n24), .Z(n387) );
  AOI22CDNM1P U94 ( .A(n24), .B(n154), .C(\Queue[4][3] ), .D(n24), .Z(n388) );
  AOI22CDNM1P U95 ( .A(n24), .B(n156), .C(\Queue[4][4] ), .D(n24), .Z(n389) );
  AOI22CDNM1P U96 ( .A(n24), .B(n158), .C(\Queue[4][5] ), .D(n24), .Z(n390) );
  AOI22CDNM1P U97 ( .A(n24), .B(n160), .C(\Queue[4][6] ), .D(n24), .Z(n391) );
  AOI22CDNM1P U98 ( .A(n24), .B(n162), .C(\Queue[4][7] ), .D(n24), .Z(n392) );
  AOI22CDNM1P U99 ( .A(n24), .B(n164), .C(\Queue[4][8] ), .D(n24), .Z(n393) );
  AOI22CDNM1P U100 ( .A(n24), .B(n166), .C(\Queue[4][9] ), .D(n24), .Z(n394)
         );
  AOI22CDNM1P U101 ( .A(n24), .B(n168), .C(\Queue[4][10] ), .D(n24), .Z(n395)
         );
  AOI22CDNM1P U102 ( .A(n24), .B(n170), .C(\Queue[4][11] ), .D(n24), .Z(n396)
         );
  AOI22CDNM1P U103 ( .A(n24), .B(n172), .C(\Queue[4][12] ), .D(n24), .Z(n397)
         );
  AOI22CDNM1P U104 ( .A(n24), .B(n174), .C(\Queue[4][13] ), .D(n24), .Z(n398)
         );
  AOI22CDNM1P U105 ( .A(n24), .B(n176), .C(\Queue[4][14] ), .D(n24), .Z(n399)
         );
  AOI22CDNM1P U106 ( .A(n24), .B(n178), .C(\Queue[4][15] ), .D(n24), .Z(n400)
         );
  AOI22CDNM1P U107 ( .A(n24), .B(n180), .C(\Queue[4][16] ), .D(n24), .Z(n401)
         );
  AOI22CDNM1P U108 ( .A(n24), .B(n182), .C(\Queue[4][17] ), .D(n24), .Z(n402)
         );
  AOI22CDNM1P U109 ( .A(n24), .B(n184), .C(\Queue[4][18] ), .D(n24), .Z(n403)
         );
  AOI22CDNM1P U110 ( .A(n24), .B(n186), .C(\Queue[4][19] ), .D(n24), .Z(n404)
         );
  AOI22CDNM1P U111 ( .A(n24), .B(n188), .C(\Queue[4][20] ), .D(n24), .Z(n405)
         );
  AOI22CDNM1P U112 ( .A(n24), .B(n190), .C(\Queue[4][21] ), .D(n24), .Z(n406)
         );
  AOI22CDNM1P U113 ( .A(n24), .B(n192), .C(\Queue[4][22] ), .D(n24), .Z(n407)
         );
  AOI22CDNM1P U114 ( .A(n24), .B(n194), .C(\Queue[4][23] ), .D(n24), .Z(n408)
         );
  AOI22CDNM1P U115 ( .A(n24), .B(n196), .C(\Queue[4][24] ), .D(n24), .Z(n409)
         );
  AOI22CDNM1P U116 ( .A(n24), .B(n198), .C(\Queue[4][25] ), .D(n24), .Z(n410)
         );
  AOI22CDNM1P U117 ( .A(n24), .B(n200), .C(\Queue[4][26] ), .D(n24), .Z(n411)
         );
  AOI22CDNM1P U118 ( .A(n24), .B(n202), .C(\Queue[4][27] ), .D(n24), .Z(n412)
         );
  AOI22CDNM1P U119 ( .A(n24), .B(n204), .C(\Queue[4][28] ), .D(n24), .Z(n413)
         );
  AOI22CDNM1P U120 ( .A(n24), .B(n206), .C(\Queue[4][29] ), .D(n24), .Z(n414)
         );
  AOI22CDNM1P U121 ( .A(n24), .B(n208), .C(\Queue[4][30] ), .D(n24), .Z(n415)
         );
  OAI22CDNM1P U122 ( .A(n143), .B(n25), .C(n378), .D(Full), .Z(n416) );
  AOI22M1P U123 ( .A(\Queue[2][0] ), .B(n7), .C(\Queue[1][0] ), .D(n4), .Z(n29) );
  OAI21M1P U124 ( .A(n148), .B(n9), .C(n29), .Z(n417) );
  AOI22M1P U125 ( .A(n6), .B(\Queue[2][1] ), .C(\Queue[1][1] ), .D(n4), .Z(n30) );
  OAI21M1P U126 ( .A(n8), .B(n150), .C(n30), .Z(n418) );
  AOI22M1P U127 ( .A(n7), .B(\Queue[2][2] ), .C(\Queue[1][2] ), .D(n4), .Z(n31) );
  OAI21M1P U128 ( .A(n9), .B(n152), .C(n31), .Z(n419) );
  AOI22M1P U129 ( .A(n7), .B(\Queue[2][3] ), .C(\Queue[1][3] ), .D(n4), .Z(n32) );
  OAI21M1P U130 ( .A(n9), .B(n154), .C(n32), .Z(n420) );
  AOI22M1P U131 ( .A(n7), .B(\Queue[2][4] ), .C(\Queue[1][4] ), .D(n4), .Z(n33) );
  OAI21M1P U132 ( .A(n9), .B(n156), .C(n33), .Z(n421) );
  AOI22M1P U133 ( .A(n7), .B(\Queue[2][5] ), .C(\Queue[1][5] ), .D(n4), .Z(n34) );
  OAI21M1P U134 ( .A(n9), .B(n158), .C(n34), .Z(n422) );
  AOI22M1P U135 ( .A(n7), .B(\Queue[2][6] ), .C(\Queue[1][6] ), .D(n4), .Z(n35) );
  OAI21M1P U136 ( .A(n9), .B(n160), .C(n35), .Z(n423) );
  AOI22M1P U137 ( .A(n7), .B(\Queue[2][7] ), .C(\Queue[1][7] ), .D(n4), .Z(n36) );
  OAI21M1P U138 ( .A(n9), .B(n162), .C(n36), .Z(n424) );
  AOI22M1P U139 ( .A(n7), .B(\Queue[2][8] ), .C(\Queue[1][8] ), .D(n4), .Z(n37) );
  OAI21M1P U140 ( .A(n9), .B(n164), .C(n37), .Z(n425) );
  AOI22M1P U141 ( .A(n7), .B(\Queue[2][9] ), .C(\Queue[1][9] ), .D(n4), .Z(n38) );
  OAI21M1P U142 ( .A(n9), .B(n166), .C(n38), .Z(n426) );
  AOI22M1P U143 ( .A(n7), .B(\Queue[2][10] ), .C(\Queue[1][10] ), .D(n5), .Z(
        n39) );
  OAI21M1P U144 ( .A(n9), .B(n168), .C(n39), .Z(n427) );
  AOI22M1P U145 ( .A(n7), .B(\Queue[2][11] ), .C(\Queue[1][11] ), .D(n4), .Z(
        n40) );
  OAI21M1P U146 ( .A(n9), .B(n170), .C(n40), .Z(n428) );
  AOI22M1P U147 ( .A(n6), .B(\Queue[2][12] ), .C(\Queue[1][12] ), .D(n60), .Z(
        n41) );
  OAI21M1P U148 ( .A(n8), .B(n172), .C(n41), .Z(n429) );
  AOI22M1P U149 ( .A(n6), .B(\Queue[2][13] ), .C(\Queue[1][13] ), .D(n60), .Z(
        n42) );
  OAI21M1P U150 ( .A(n8), .B(n174), .C(n42), .Z(n430) );
  AOI22M1P U151 ( .A(n6), .B(\Queue[2][14] ), .C(\Queue[1][14] ), .D(n60), .Z(
        n43) );
  OAI21M1P U152 ( .A(n8), .B(n176), .C(n43), .Z(n431) );
  AOI22M1P U153 ( .A(n6), .B(\Queue[2][15] ), .C(\Queue[1][15] ), .D(n60), .Z(
        n44) );
  OAI21M1P U154 ( .A(n8), .B(n178), .C(n44), .Z(n432) );
  AOI22M1P U155 ( .A(n6), .B(\Queue[2][16] ), .C(\Queue[1][16] ), .D(n60), .Z(
        n45) );
  OAI21M1P U156 ( .A(n8), .B(n180), .C(n45), .Z(n433) );
  AOI22M1P U157 ( .A(n6), .B(\Queue[2][17] ), .C(\Queue[1][17] ), .D(n60), .Z(
        n46) );
  OAI21M1P U158 ( .A(n8), .B(n182), .C(n46), .Z(n434) );
  AOI22M1P U159 ( .A(n6), .B(\Queue[2][18] ), .C(\Queue[1][18] ), .D(n5), .Z(
        n47) );
  OAI21M1P U160 ( .A(n8), .B(n184), .C(n47), .Z(n435) );
  AOI22M1P U161 ( .A(n6), .B(\Queue[2][19] ), .C(\Queue[1][19] ), .D(n5), .Z(
        n48) );
  OAI21M1P U162 ( .A(n8), .B(n186), .C(n48), .Z(n436) );
  AOI22M1P U163 ( .A(n6), .B(\Queue[2][20] ), .C(\Queue[1][20] ), .D(n5), .Z(
        n49) );
  OAI21M1P U164 ( .A(n8), .B(n188), .C(n49), .Z(n437) );
  AOI22M1P U165 ( .A(n6), .B(\Queue[2][21] ), .C(\Queue[1][21] ), .D(n5), .Z(
        n50) );
  OAI21M1P U166 ( .A(n8), .B(n190), .C(n50), .Z(n438) );
  AOI22M1P U167 ( .A(n7), .B(\Queue[2][22] ), .C(\Queue[1][22] ), .D(n5), .Z(
        n51) );
  OAI21M1P U168 ( .A(n8), .B(n192), .C(n51), .Z(n439) );
  AOI22M1P U169 ( .A(n6), .B(\Queue[2][23] ), .C(\Queue[1][23] ), .D(n5), .Z(
        n52) );
  OAI21M1P U170 ( .A(n8), .B(n194), .C(n52), .Z(n440) );
  AOI22M1P U171 ( .A(n7), .B(\Queue[2][24] ), .C(\Queue[1][24] ), .D(n5), .Z(
        n53) );
  OAI21M1P U172 ( .A(n8), .B(n196), .C(n53), .Z(n441) );
  AOI22M1P U173 ( .A(n61), .B(\Queue[2][25] ), .C(\Queue[1][25] ), .D(n5), .Z(
        n54) );
  OAI21M1P U174 ( .A(n8), .B(n198), .C(n54), .Z(n442) );
  AOI22M1P U175 ( .A(n61), .B(\Queue[2][26] ), .C(\Queue[1][26] ), .D(n5), .Z(
        n55) );
  OAI21M1P U176 ( .A(n8), .B(n200), .C(n55), .Z(n443) );
  AOI22M1P U177 ( .A(n61), .B(\Queue[2][27] ), .C(\Queue[1][27] ), .D(n5), .Z(
        n56) );
  OAI21M1P U178 ( .A(n8), .B(n202), .C(n56), .Z(n444) );
  AOI22M1P U179 ( .A(n61), .B(\Queue[2][28] ), .C(\Queue[1][28] ), .D(n4), .Z(
        n57) );
  OAI21M1P U180 ( .A(n8), .B(n204), .C(n57), .Z(n445) );
  AOI22M1P U181 ( .A(n61), .B(\Queue[2][29] ), .C(\Queue[1][29] ), .D(n60), 
        .Z(n58) );
  OAI21M1P U182 ( .A(n8), .B(n206), .C(n58), .Z(n446) );
  AOI22M1P U183 ( .A(n61), .B(\Queue[2][30] ), .C(\Queue[1][30] ), .D(n5), .Z(
        n59) );
  OAI21M1P U184 ( .A(n8), .B(n208), .C(n59), .Z(n447) );
  AOI22M1P U185 ( .A(n61), .B(\Queue[2][31] ), .C(\Queue[1][31] ), .D(n4), .Z(
        n62) );
  OAI21M1P U186 ( .A(n8), .B(n377), .C(n62), .Z(n448) );
  AOI22M1P U187 ( .A(\Queue[1][0] ), .B(n99), .C(n98), .D(Packet_Out[0]), .Z(
        n67) );
  OAI21M1P U188 ( .A(n148), .B(n10), .C(n67), .Z(n449) );
  AOI22M1P U189 ( .A(\Queue[1][1] ), .B(n99), .C(n98), .D(Packet_Out[1]), .Z(
        n68) );
  OAI21M1P U190 ( .A(n150), .B(n10), .C(n68), .Z(n450) );
  AOI22M1P U191 ( .A(\Queue[1][2] ), .B(n99), .C(n98), .D(Packet_Out[2]), .Z(
        n69) );
  OAI21M1P U192 ( .A(n152), .B(n10), .C(n69), .Z(n451) );
  AOI22M1P U193 ( .A(\Queue[1][3] ), .B(n99), .C(n98), .D(Packet_Out[3]), .Z(
        n70) );
  OAI21M1P U194 ( .A(n154), .B(n10), .C(n70), .Z(n452) );
  AOI22M1P U195 ( .A(\Queue[1][4] ), .B(n99), .C(n98), .D(Packet_Out[4]), .Z(
        n71) );
  OAI21M1P U196 ( .A(n156), .B(n10), .C(n71), .Z(n453) );
  AOI22M1P U197 ( .A(\Queue[1][5] ), .B(n99), .C(n98), .D(Packet_Out[5]), .Z(
        n72) );
  OAI21M1P U198 ( .A(n158), .B(n10), .C(n72), .Z(n454) );
  AOI22M1P U199 ( .A(\Queue[1][6] ), .B(n99), .C(n98), .D(Packet_Out[6]), .Z(
        n73) );
  OAI21M1P U200 ( .A(n160), .B(n10), .C(n73), .Z(n455) );
  AOI22M1P U201 ( .A(\Queue[1][7] ), .B(n99), .C(n98), .D(Packet_Out[7]), .Z(
        n74) );
  OAI21M1P U202 ( .A(n162), .B(n10), .C(n74), .Z(n456) );
  AOI22M1P U203 ( .A(\Queue[1][8] ), .B(n99), .C(n98), .D(Packet_Out[8]), .Z(
        n75) );
  OAI21M1P U204 ( .A(n164), .B(n10), .C(n75), .Z(n457) );
  AOI22M1P U205 ( .A(\Queue[1][9] ), .B(n99), .C(n98), .D(Packet_Out[9]), .Z(
        n76) );
  OAI21M1P U206 ( .A(n166), .B(n10), .C(n76), .Z(n458) );
  AOI22M1P U207 ( .A(\Queue[1][10] ), .B(n99), .C(n98), .D(Packet_Out[10]), 
        .Z(n77) );
  OAI21M1P U208 ( .A(n168), .B(n10), .C(n77), .Z(n459) );
  AOI22M1P U209 ( .A(\Queue[1][11] ), .B(n99), .C(n98), .D(Packet_Out[11]), 
        .Z(n78) );
  OAI21M1P U210 ( .A(n170), .B(n10), .C(n78), .Z(n460) );
  AOI22M1P U211 ( .A(\Queue[1][12] ), .B(n99), .C(n98), .D(Packet_Out[12]), 
        .Z(n79) );
  OAI21M1P U212 ( .A(n172), .B(n10), .C(n79), .Z(n461) );
  AOI22M1P U213 ( .A(\Queue[1][13] ), .B(n99), .C(n98), .D(Packet_Out[13]), 
        .Z(n80) );
  OAI21M1P U214 ( .A(n174), .B(n10), .C(n80), .Z(n462) );
  AOI22M1P U215 ( .A(\Queue[1][14] ), .B(n99), .C(n98), .D(Packet_Out[14]), 
        .Z(n81) );
  OAI21M1P U216 ( .A(n176), .B(n10), .C(n81), .Z(n463) );
  AOI22M1P U217 ( .A(\Queue[1][15] ), .B(n99), .C(n98), .D(Packet_Out[15]), 
        .Z(n82) );
  OAI21M1P U218 ( .A(n178), .B(n10), .C(n82), .Z(n464) );
  AOI22M1P U219 ( .A(\Queue[1][16] ), .B(n99), .C(n98), .D(Packet_Out[16]), 
        .Z(n83) );
  OAI21M1P U220 ( .A(n180), .B(n10), .C(n83), .Z(n465) );
  AOI22M1P U221 ( .A(\Queue[1][17] ), .B(n99), .C(n98), .D(Packet_Out[17]), 
        .Z(n84) );
  OAI21M1P U222 ( .A(n182), .B(n10), .C(n84), .Z(n466) );
  AOI22M1P U223 ( .A(\Queue[1][18] ), .B(n99), .C(n98), .D(Packet_Out[18]), 
        .Z(n85) );
  OAI21M1P U224 ( .A(n184), .B(n10), .C(n85), .Z(n467) );
  AOI22M1P U225 ( .A(\Queue[1][19] ), .B(n99), .C(n98), .D(Packet_Out[19]), 
        .Z(n86) );
  OAI21M1P U226 ( .A(n186), .B(n10), .C(n86), .Z(n468) );
  AOI22M1P U227 ( .A(\Queue[1][20] ), .B(n99), .C(n98), .D(Packet_Out[20]), 
        .Z(n87) );
  OAI21M1P U228 ( .A(n188), .B(n11), .C(n87), .Z(n469) );
  AOI22M1P U229 ( .A(\Queue[1][21] ), .B(n99), .C(n98), .D(Packet_Out[21]), 
        .Z(n88) );
  OAI21M1P U230 ( .A(n190), .B(n11), .C(n88), .Z(n470) );
  AOI22M1P U231 ( .A(\Queue[1][22] ), .B(n99), .C(n98), .D(Packet_Out[22]), 
        .Z(n89) );
  OAI21M1P U232 ( .A(n192), .B(n11), .C(n89), .Z(n471) );
  AOI22M1P U233 ( .A(\Queue[1][23] ), .B(n99), .C(n98), .D(Packet_Out[23]), 
        .Z(n90) );
  OAI21M1P U234 ( .A(n194), .B(n11), .C(n90), .Z(n472) );
  AOI22M1P U235 ( .A(\Queue[1][24] ), .B(n99), .C(n98), .D(Packet_Out[24]), 
        .Z(n91) );
  OAI21M1P U236 ( .A(n196), .B(n11), .C(n91), .Z(n473) );
  AOI22M1P U237 ( .A(\Queue[1][25] ), .B(n99), .C(n98), .D(Packet_Out[25]), 
        .Z(n92) );
  OAI21M1P U238 ( .A(n198), .B(n11), .C(n92), .Z(n474) );
  AOI22M1P U239 ( .A(\Queue[1][26] ), .B(n99), .C(n98), .D(Packet_Out[26]), 
        .Z(n93) );
  OAI21M1P U240 ( .A(n200), .B(n11), .C(n93), .Z(n475) );
  AOI22M1P U241 ( .A(\Queue[1][27] ), .B(n99), .C(n98), .D(Packet_Out[27]), 
        .Z(n94) );
  OAI21M1P U242 ( .A(n202), .B(n11), .C(n94), .Z(n476) );
  AOI22M1P U243 ( .A(\Queue[1][28] ), .B(n99), .C(n98), .D(Packet_Out[28]), 
        .Z(n95) );
  OAI21M1P U244 ( .A(n204), .B(n11), .C(n95), .Z(n477) );
  AOI22M1P U245 ( .A(\Queue[1][29] ), .B(n99), .C(n98), .D(Packet_Out[29]), 
        .Z(n96) );
  OAI21M1P U246 ( .A(n206), .B(n11), .C(n96), .Z(n478) );
  AOI22M1P U247 ( .A(\Queue[1][30] ), .B(n99), .C(n98), .D(Packet_Out[30]), 
        .Z(n97) );
  OAI21M1P U248 ( .A(n208), .B(n11), .C(n97), .Z(n479) );
  AOI22M1P U249 ( .A(\Queue[1][31] ), .B(n99), .C(n98), .D(Packet_Out[31]), 
        .Z(n100) );
  OAI21M1P U250 ( .A(n377), .B(n10), .C(n100), .Z(n480) );
  ND2M1P U251 ( .A(n103), .B(n141), .Z(n142) );
  AOI21M1P U252 ( .A(Write_Ack), .B(n144), .C(n145), .Z(n136) );
  AOI22M1P U253 ( .A(\Queue[2][0] ), .B(n13), .C(\Queue[3][0] ), .D(n12), .Z(
        n105) );
  OAI21M1P U254 ( .A(n148), .B(n139), .C(n105), .Z(n481) );
  AOI22M1P U255 ( .A(\Queue[2][1] ), .B(n13), .C(n3), .D(\Queue[3][1] ), .Z(
        n106) );
  OAI21M1P U256 ( .A(n150), .B(n139), .C(n106), .Z(n482) );
  AOI22M1P U257 ( .A(\Queue[2][2] ), .B(n13), .C(n12), .D(\Queue[3][2] ), .Z(
        n107) );
  OAI21M1P U258 ( .A(n152), .B(n139), .C(n107), .Z(n483) );
  AOI22M1P U259 ( .A(\Queue[2][3] ), .B(n13), .C(n12), .D(\Queue[3][3] ), .Z(
        n108) );
  OAI21M1P U260 ( .A(n154), .B(n139), .C(n108), .Z(n484) );
  AOI22M1P U261 ( .A(\Queue[2][4] ), .B(n13), .C(n12), .D(\Queue[3][4] ), .Z(
        n109) );
  OAI21M1P U262 ( .A(n156), .B(n139), .C(n109), .Z(n485) );
  AOI22M1P U263 ( .A(\Queue[2][5] ), .B(n13), .C(n12), .D(\Queue[3][5] ), .Z(
        n110) );
  OAI21M1P U264 ( .A(n158), .B(n139), .C(n110), .Z(n486) );
  AOI22M1P U265 ( .A(\Queue[2][6] ), .B(n13), .C(n12), .D(\Queue[3][6] ), .Z(
        n111) );
  OAI21M1P U266 ( .A(n160), .B(n139), .C(n111), .Z(n487) );
  AOI22M1P U267 ( .A(\Queue[2][7] ), .B(n13), .C(n12), .D(\Queue[3][7] ), .Z(
        n112) );
  OAI21M1P U268 ( .A(n162), .B(n139), .C(n112), .Z(n488) );
  AOI22M1P U269 ( .A(\Queue[2][8] ), .B(n13), .C(n12), .D(\Queue[3][8] ), .Z(
        n113) );
  OAI21M1P U270 ( .A(n164), .B(n139), .C(n113), .Z(n489) );
  AOI22M1P U271 ( .A(\Queue[2][9] ), .B(n13), .C(n12), .D(\Queue[3][9] ), .Z(
        n114) );
  OAI21M1P U272 ( .A(n166), .B(n139), .C(n114), .Z(n490) );
  AOI22M1P U273 ( .A(\Queue[2][10] ), .B(n13), .C(n12), .D(\Queue[3][10] ), 
        .Z(n115) );
  OAI21M1P U274 ( .A(n168), .B(n139), .C(n115), .Z(n491) );
  AOI22M1P U275 ( .A(\Queue[2][11] ), .B(n13), .C(n12), .D(\Queue[3][11] ), 
        .Z(n116) );
  OAI21M1P U276 ( .A(n170), .B(n139), .C(n116), .Z(n492) );
  AOI22M1P U277 ( .A(\Queue[2][12] ), .B(n13), .C(n3), .D(\Queue[3][12] ), .Z(
        n117) );
  OAI21M1P U278 ( .A(n172), .B(n139), .C(n117), .Z(n493) );
  AOI22M1P U279 ( .A(\Queue[2][13] ), .B(n13), .C(n3), .D(\Queue[3][13] ), .Z(
        n118) );
  OAI21M1P U280 ( .A(n174), .B(n139), .C(n118), .Z(n494) );
  AOI22M1P U281 ( .A(\Queue[2][14] ), .B(n13), .C(n3), .D(\Queue[3][14] ), .Z(
        n119) );
  OAI21M1P U282 ( .A(n176), .B(n139), .C(n119), .Z(n495) );
  AOI22M1P U283 ( .A(\Queue[2][15] ), .B(n13), .C(n3), .D(\Queue[3][15] ), .Z(
        n120) );
  OAI21M1P U284 ( .A(n178), .B(n139), .C(n120), .Z(n496) );
  AOI22M1P U285 ( .A(\Queue[2][16] ), .B(n13), .C(n3), .D(\Queue[3][16] ), .Z(
        n121) );
  OAI21M1P U286 ( .A(n180), .B(n139), .C(n121), .Z(n497) );
  AOI22M1P U287 ( .A(\Queue[2][17] ), .B(n13), .C(n3), .D(\Queue[3][17] ), .Z(
        n122) );
  OAI21M1P U288 ( .A(n182), .B(n139), .C(n122), .Z(n498) );
  AOI22M1P U289 ( .A(\Queue[2][18] ), .B(n13), .C(n3), .D(\Queue[3][18] ), .Z(
        n123) );
  OAI21M1P U290 ( .A(n184), .B(n139), .C(n123), .Z(n499) );
  AOI22M1P U291 ( .A(\Queue[2][19] ), .B(n13), .C(n3), .D(\Queue[3][19] ), .Z(
        n124) );
  OAI21M1P U292 ( .A(n186), .B(n139), .C(n124), .Z(n500) );
  AOI22M1P U293 ( .A(\Queue[2][20] ), .B(n14), .C(n3), .D(\Queue[3][20] ), .Z(
        n125) );
  OAI21M1P U294 ( .A(n188), .B(n139), .C(n125), .Z(n501) );
  AOI22M1P U295 ( .A(\Queue[2][21] ), .B(n14), .C(n3), .D(\Queue[3][21] ), .Z(
        n126) );
  OAI21M1P U296 ( .A(n190), .B(n139), .C(n126), .Z(n502) );
  AOI22M1P U297 ( .A(\Queue[2][22] ), .B(n14), .C(n3), .D(\Queue[3][22] ), .Z(
        n127) );
  OAI21M1P U298 ( .A(n192), .B(n139), .C(n127), .Z(n503) );
  AOI22M1P U299 ( .A(\Queue[2][23] ), .B(n14), .C(n3), .D(\Queue[3][23] ), .Z(
        n128) );
  OAI21M1P U300 ( .A(n194), .B(n139), .C(n128), .Z(n504) );
  AOI22M1P U301 ( .A(\Queue[2][24] ), .B(n14), .C(n3), .D(\Queue[3][24] ), .Z(
        n129) );
  OAI21M1P U302 ( .A(n196), .B(n139), .C(n129), .Z(n505) );
  AOI22M1P U303 ( .A(\Queue[2][25] ), .B(n14), .C(n3), .D(\Queue[3][25] ), .Z(
        n130) );
  OAI21M1P U304 ( .A(n198), .B(n139), .C(n130), .Z(n506) );
  AOI22M1P U305 ( .A(\Queue[2][26] ), .B(n14), .C(n3), .D(\Queue[3][26] ), .Z(
        n131) );
  OAI21M1P U306 ( .A(n200), .B(n139), .C(n131), .Z(n507) );
  AOI22M1P U307 ( .A(\Queue[2][27] ), .B(n14), .C(n3), .D(\Queue[3][27] ), .Z(
        n132) );
  OAI21M1P U308 ( .A(n202), .B(n139), .C(n132), .Z(n508) );
  AOI22M1P U309 ( .A(\Queue[2][28] ), .B(n14), .C(n3), .D(\Queue[3][28] ), .Z(
        n133) );
  OAI21M1P U310 ( .A(n204), .B(n139), .C(n133), .Z(n509) );
  AOI22M1P U311 ( .A(\Queue[2][29] ), .B(n14), .C(n3), .D(\Queue[3][29] ), .Z(
        n134) );
  OAI21M1P U312 ( .A(n206), .B(n139), .C(n134), .Z(n510) );
  AOI22M1P U313 ( .A(\Queue[2][30] ), .B(n13), .C(n3), .D(\Queue[3][30] ), .Z(
        n135) );
  OAI21M1P U314 ( .A(n208), .B(n139), .C(n135), .Z(n511) );
  AOI22M1P U315 ( .A(\Queue[2][31] ), .B(n14), .C(n3), .D(\Queue[3][31] ), .Z(
        n138) );
  OAI21M1P U316 ( .A(n377), .B(n139), .C(n138), .Z(n512) );
  AOI22M1P U317 ( .A(\Queue[3][0] ), .B(n15), .C(n373), .D(\Queue[4][0] ), .Z(
        n147) );
  OAI21M1P U318 ( .A(n148), .B(n376), .C(n147), .Z(n513) );
  AOI22M1P U319 ( .A(\Queue[3][1] ), .B(n15), .C(n373), .D(\Queue[4][1] ), .Z(
        n149) );
  OAI21M1P U320 ( .A(n150), .B(n376), .C(n149), .Z(n514) );
  AOI22M1P U321 ( .A(\Queue[3][2] ), .B(n15), .C(n373), .D(\Queue[4][2] ), .Z(
        n151) );
  OAI21M1P U322 ( .A(n152), .B(n376), .C(n151), .Z(n515) );
  AOI22M1P U323 ( .A(\Queue[3][3] ), .B(n15), .C(n373), .D(\Queue[4][3] ), .Z(
        n153) );
  OAI21M1P U324 ( .A(n154), .B(n376), .C(n153), .Z(n516) );
  AOI22M1P U325 ( .A(\Queue[3][4] ), .B(n15), .C(n373), .D(\Queue[4][4] ), .Z(
        n155) );
  OAI21M1P U326 ( .A(n156), .B(n376), .C(n155), .Z(n517) );
  AOI22M1P U327 ( .A(\Queue[3][5] ), .B(n15), .C(n373), .D(\Queue[4][5] ), .Z(
        n157) );
  OAI21M1P U328 ( .A(n158), .B(n376), .C(n157), .Z(n518) );
  AOI22M1P U329 ( .A(\Queue[3][6] ), .B(n15), .C(n373), .D(\Queue[4][6] ), .Z(
        n159) );
  OAI21M1P U330 ( .A(n160), .B(n376), .C(n159), .Z(n519) );
  AOI22M1P U331 ( .A(\Queue[3][7] ), .B(n15), .C(n373), .D(\Queue[4][7] ), .Z(
        n161) );
  OAI21M1P U332 ( .A(n162), .B(n376), .C(n161), .Z(n520) );
  AOI22M1P U333 ( .A(\Queue[3][8] ), .B(n15), .C(n373), .D(\Queue[4][8] ), .Z(
        n163) );
  OAI21M1P U334 ( .A(n164), .B(n376), .C(n163), .Z(n521) );
  AOI22M1P U335 ( .A(\Queue[3][9] ), .B(n15), .C(n373), .D(\Queue[4][9] ), .Z(
        n165) );
  OAI21M1P U336 ( .A(n166), .B(n376), .C(n165), .Z(n522) );
  AOI22M1P U337 ( .A(\Queue[3][10] ), .B(n15), .C(n373), .D(\Queue[4][10] ), 
        .Z(n167) );
  OAI21M1P U338 ( .A(n168), .B(n376), .C(n167), .Z(n523) );
  AOI22M1P U339 ( .A(\Queue[3][11] ), .B(n15), .C(n373), .D(\Queue[4][11] ), 
        .Z(n169) );
  OAI21M1P U340 ( .A(n170), .B(n376), .C(n169), .Z(n524) );
  AOI22M1P U341 ( .A(\Queue[3][12] ), .B(n15), .C(n373), .D(\Queue[4][12] ), 
        .Z(n171) );
  OAI21M1P U342 ( .A(n172), .B(n376), .C(n171), .Z(n525) );
  AOI22M1P U343 ( .A(\Queue[3][13] ), .B(n15), .C(n373), .D(\Queue[4][13] ), 
        .Z(n173) );
  OAI21M1P U344 ( .A(n174), .B(n376), .C(n173), .Z(n526) );
  AOI22M1P U345 ( .A(\Queue[3][14] ), .B(n15), .C(n373), .D(\Queue[4][14] ), 
        .Z(n175) );
  OAI21M1P U346 ( .A(n176), .B(n376), .C(n175), .Z(n527) );
  AOI22M1P U347 ( .A(\Queue[3][15] ), .B(n15), .C(n373), .D(\Queue[4][15] ), 
        .Z(n177) );
  OAI21M1P U348 ( .A(n178), .B(n376), .C(n177), .Z(n528) );
  AOI22M1P U349 ( .A(\Queue[3][16] ), .B(n15), .C(n373), .D(\Queue[4][16] ), 
        .Z(n179) );
  OAI21M1P U350 ( .A(n180), .B(n376), .C(n179), .Z(n529) );
  AOI22M1P U351 ( .A(\Queue[3][17] ), .B(n15), .C(n373), .D(\Queue[4][17] ), 
        .Z(n181) );
  OAI21M1P U352 ( .A(n182), .B(n376), .C(n181), .Z(n530) );
  AOI22M1P U353 ( .A(\Queue[3][18] ), .B(n15), .C(n373), .D(\Queue[4][18] ), 
        .Z(n183) );
  OAI21M1P U354 ( .A(n184), .B(n376), .C(n183), .Z(n531) );
  AOI22M1P U355 ( .A(\Queue[3][19] ), .B(n15), .C(n373), .D(\Queue[4][19] ), 
        .Z(n185) );
  OAI21M1P U356 ( .A(n186), .B(n376), .C(n185), .Z(n532) );
  AOI22M1P U357 ( .A(\Queue[3][20] ), .B(n16), .C(n373), .D(\Queue[4][20] ), 
        .Z(n187) );
  OAI21M1P U358 ( .A(n188), .B(n376), .C(n187), .Z(n533) );
  AOI22M1P U359 ( .A(\Queue[3][21] ), .B(n16), .C(n373), .D(\Queue[4][21] ), 
        .Z(n189) );
  OAI21M1P U360 ( .A(n190), .B(n376), .C(n189), .Z(n534) );
  AOI22M1P U361 ( .A(\Queue[3][22] ), .B(n16), .C(n373), .D(\Queue[4][22] ), 
        .Z(n191) );
  OAI21M1P U362 ( .A(n192), .B(n376), .C(n191), .Z(n535) );
  AOI22M1P U363 ( .A(\Queue[3][23] ), .B(n16), .C(n373), .D(\Queue[4][23] ), 
        .Z(n193) );
  OAI21M1P U364 ( .A(n194), .B(n376), .C(n193), .Z(n536) );
  AOI22M1P U365 ( .A(\Queue[3][24] ), .B(n16), .C(n373), .D(\Queue[4][24] ), 
        .Z(n195) );
  OAI21M1P U366 ( .A(n196), .B(n376), .C(n195), .Z(n537) );
  AOI22M1P U367 ( .A(\Queue[3][25] ), .B(n16), .C(n373), .D(\Queue[4][25] ), 
        .Z(n197) );
  OAI21M1P U368 ( .A(n198), .B(n376), .C(n197), .Z(n538) );
  AOI22M1P U369 ( .A(\Queue[3][26] ), .B(n16), .C(n373), .D(\Queue[4][26] ), 
        .Z(n199) );
  OAI21M1P U370 ( .A(n200), .B(n376), .C(n199), .Z(n539) );
  AOI22M1P U371 ( .A(\Queue[3][27] ), .B(n16), .C(n373), .D(\Queue[4][27] ), 
        .Z(n201) );
  OAI21M1P U372 ( .A(n202), .B(n376), .C(n201), .Z(n540) );
  AOI22M1P U373 ( .A(\Queue[3][28] ), .B(n16), .C(n373), .D(\Queue[4][28] ), 
        .Z(n203) );
  OAI21M1P U374 ( .A(n204), .B(n376), .C(n203), .Z(n541) );
  AOI22M1P U375 ( .A(\Queue[3][29] ), .B(n16), .C(n373), .D(\Queue[4][29] ), 
        .Z(n205) );
  OAI21M1P U376 ( .A(n206), .B(n376), .C(n205), .Z(n542) );
  AOI22M1P U377 ( .A(\Queue[3][30] ), .B(n15), .C(n373), .D(\Queue[4][30] ), 
        .Z(n207) );
  OAI21M1P U378 ( .A(n208), .B(n376), .C(n207), .Z(n543) );
  AOI22M1P U379 ( .A(\Queue[3][31] ), .B(n16), .C(n373), .D(\Queue[4][31] ), 
        .Z(n375) );
  OAI21M1P U380 ( .A(n377), .B(n376), .C(n375), .Z(n544) );
  N1M1P U381 ( .A(n545), .Z(Empty) );
  AOI22M1P U382 ( .A(n380), .B(n379), .C(n378), .D(Empty), .Z(n546) );
endmodule


module Link_Control_0 ( Clk_r, Rst_n, Tx_Ready, Tx_Error, RxData_Valid, RxData, 
        Packet_From_Core, TxQueue_Write, RxQueue_Read, TxData_Valid, TxData, 
        Error_Ack, Core_Rcv_Ready, Packet_To_Core, RxQueue_Empty, TxQueue_Full
 );
  input [31:0] RxData;
  input [31:0] Packet_From_Core;
  output [31:0] TxData;
  output [31:0] Packet_To_Core;
  input Clk_r, Rst_n, Tx_Ready, Tx_Error, RxData_Valid, TxQueue_Write,
         RxQueue_Read;
  output TxData_Valid, Error_Ack, Core_Rcv_Ready, RxQueue_Empty, TxQueue_Full;
  wire   TxQueue_Read, TxQueue_Empty, RxQueue_Write, RxQueue_Full, N9, N16, n1,
         n2, n3, n4, n5;

  Packet_Queue_0 TxQueue ( .Clk_r(Clk_r), .Rst_n(Rst_n), .Packet_In(
        Packet_From_Core), .Read_Ack(TxQueue_Read), .Write_Ack(TxQueue_Write), 
        .Packet_Out(TxData), .Empty(TxQueue_Empty), .Full(TxQueue_Full) );
  Packet_Queue_9 RxQueue ( .Clk_r(Clk_r), .Rst_n(Rst_n), .Packet_In(RxData), 
        .Read_Ack(RxQueue_Read), .Write_Ack(RxQueue_Write), .Packet_Out(
        Packet_To_Core), .Empty(RxQueue_Empty), .Full(RxQueue_Full) );
  FD4QM1P TxData_Valid_reg ( .D(n1), .CP(Clk_r), .SD(Rst_n), .Q(n2) );
  FD2QM1P Error_Ack_reg ( .D(Tx_Error), .CP(Clk_r), .CD(Rst_n), .Q(Error_Ack)
         );
  FD4QM1P RxQueue_Write_reg ( .D(n3), .CP(Clk_r), .SD(Rst_n), .Q(n4) );
  FD2QM1P TxQueue_Read_reg ( .D(N16), .CP(Clk_r), .CD(Rst_n), .Q(TxQueue_Read)
         );
  FD2QM1P Core_Rcv_Ready_reg ( .D(N9), .CP(Clk_r), .CD(Rst_n), .Q(
        Core_Rcv_Ready) );
  N1M3P U3 ( .A(n4), .Z(RxQueue_Write) );
  OA21M1P U4 ( .A(Core_Rcv_Ready), .B(n5), .C(n4), .Z(N9) );
  NR2M1P U5 ( .A(n2), .B(Tx_Ready), .Z(N16) );
  NR2M1P U6 ( .A(RxData_Valid), .B(RxQueue_Full), .Z(n5) );
  N1M1P U7 ( .A(n2), .Z(TxData_Valid) );
  ND3M1P U8 ( .A(n4), .B(Core_Rcv_Ready), .C(RxData_Valid), .Z(n3) );
  AO21CNM1P U9 ( .A(n2), .B(TxQueue_Empty), .C(Tx_Ready), .Z(n1) );
endmodule


module Routing_State_Machine ( Clk_r, Rst_n, Router_Address, Link_Config, 
        Packet_From_Link_N, Packet_From_Link_S, Packet_From_Link_W, 
        Packet_From_Link_E, Packet_From_Node, RxQueue_Empty_N, RxQueue_Empty_S, 
        RxQueue_Empty_W, RxQueue_Empty_E, TxQueue_Full_N, TxQueue_Full_S, 
        TxQueue_Full_W, TxQueue_Full_E, To_Node_Full, Node_Queue_Empty, 
        Packet_To_Link_N, Packet_To_Link_S, Packet_To_Link_W, Packet_To_Link_E, 
        Packet_To_Node, TxQueue_Write_N, TxQueue_Write_S, TxQueue_Write_W, 
        TxQueue_Write_E, To_Node_Write, RxQueue_Read_N, RxQueue_Read_S, 
        RxQueue_Read_W, RxQueue_Read_E, Node_Read );
  input [7:0] Router_Address;
  input [3:0] Link_Config;
  input [31:0] Packet_From_Link_N;
  input [31:0] Packet_From_Link_S;
  input [31:0] Packet_From_Link_W;
  input [31:0] Packet_From_Link_E;
  input [31:0] Packet_From_Node;
  output [31:0] Packet_To_Link_N;
  output [31:0] Packet_To_Link_S;
  output [31:0] Packet_To_Link_W;
  output [31:0] Packet_To_Link_E;
  output [31:0] Packet_To_Node;
  input Clk_r, Rst_n, RxQueue_Empty_N, RxQueue_Empty_S, RxQueue_Empty_W,
         RxQueue_Empty_E, TxQueue_Full_N, TxQueue_Full_S, TxQueue_Full_W,
         TxQueue_Full_E, To_Node_Full, Node_Queue_Empty;
  output TxQueue_Write_N, TxQueue_Write_S, TxQueue_Write_W, TxQueue_Write_E,
         To_Node_Write, RxQueue_Read_N, RxQueue_Read_S, RxQueue_Read_W,
         RxQueue_Read_E, Node_Read;
  wire   Packet_From_Node_31, Packet_From_Node_30, Packet_From_Node_29,
         Packet_From_Node_28, Packet_From_Node_27, Packet_From_Node_26,
         Packet_From_Node_25, Packet_From_Node_24, N43, N44, N48, N108, N109,
         N110, N111, N112, N113, N114, N115, n1, n2, n3, n4, n5, n6, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n32, n33, n34, n35, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n57, n107, n245, n246, n247, n249,
         n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
         n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n31, n36, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n248, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299;
  wire   [31:0] chosenPacket;
  wire   [2:0] dataLocation;
  assign Packet_From_Node_31 = Packet_From_Node[31];
  assign Packet_From_Node_30 = Packet_From_Node[30];
  assign Packet_From_Node_29 = Packet_From_Node[29];
  assign Packet_From_Node_28 = Packet_From_Node[28];
  assign Packet_From_Node_27 = Packet_From_Node[27];
  assign Packet_From_Node_26 = Packet_From_Node[26];
  assign Packet_From_Node_25 = Packet_From_Node[25];
  assign Packet_From_Node_24 = Packet_From_Node[24];

  FD2LQM1P \dataLocation_reg[0]  ( .D(N43), .LD(n8), .CP(Clk_r), .CD(Rst_n), 
        .Q(dataLocation[0]) );
  FD4QM1P \Packet_To_Node_reg[16]  ( .D(n25), .CP(Clk_r), .SD(Rst_n), .Q(
        Packet_To_Node[16]) );
  FD4QM1P \Packet_To_Node_reg[17]  ( .D(n26), .CP(Clk_r), .SD(Rst_n), .Q(
        Packet_To_Node[17]) );
  FD4QM1P \Packet_To_Node_reg[18]  ( .D(n27), .CP(Clk_r), .SD(Rst_n), .Q(
        Packet_To_Node[18]) );
  FD4QM1P \Packet_To_Node_reg[19]  ( .D(n28), .CP(Clk_r), .SD(Rst_n), .Q(
        Packet_To_Node[19]) );
  FD4QM1P \Packet_To_Node_reg[20]  ( .D(n29), .CP(Clk_r), .SD(Rst_n), .Q(
        Packet_To_Node[20]) );
  FD4QM1P \Packet_To_Node_reg[21]  ( .D(n30), .CP(Clk_r), .SD(Rst_n), .Q(
        Packet_To_Node[21]) );
  FD4QM1P \Packet_To_Node_reg[23]  ( .D(n32), .CP(Clk_r), .SD(Rst_n), .Q(
        Packet_To_Node[23]) );
  FD2LQM1P \dataLocation_reg[1]  ( .D(N44), .LD(n8), .CP(Clk_r), .CD(Rst_n), 
        .Q(dataLocation[1]) );
  FD2LQM1P \dataLocation_reg[2]  ( .D(n57), .LD(n8), .CP(Clk_r), .CD(Rst_n), 
        .Q(n6) );
  FD1QM1P \chosenPacket_reg[31]  ( .D(n263), .CP(Clk_r), .Q(chosenPacket[31])
         );
  FD2LQM1P \Packet_To_Node_reg[31]  ( .D(n41), .LD(n58), .CP(Clk_r), .CD(Rst_n), .Q(n5) );
  FD1QM1P \chosenPacket_reg[30]  ( .D(n264), .CP(Clk_r), .Q(chosenPacket[30])
         );
  FD2LQM1P \Packet_To_Node_reg[30]  ( .D(n42), .LD(n58), .CP(Clk_r), .CD(Rst_n), .Q(n4) );
  FD1QM1P \chosenPacket_reg[29]  ( .D(n265), .CP(Clk_r), .Q(chosenPacket[29])
         );
  FD2LQM1P \Packet_To_Node_reg[29]  ( .D(n43), .LD(n58), .CP(Clk_r), .CD(Rst_n), .Q(n3) );
  FD1QM1P \chosenPacket_reg[28]  ( .D(n266), .CP(Clk_r), .Q(chosenPacket[28])
         );
  FD4QM1P \Packet_To_Node_reg[28]  ( .D(n35), .CP(Clk_r), .SD(Rst_n), .Q(
        Packet_To_Node[28]) );
  FD1QM1P \chosenPacket_reg[27]  ( .D(n267), .CP(Clk_r), .Q(chosenPacket[27])
         );
  FD2LQM1P \Packet_To_Node_reg[27]  ( .D(n44), .LD(n58), .CP(Clk_r), .CD(Rst_n), .Q(n2) );
  FD1QM1P \chosenPacket_reg[26]  ( .D(n268), .CP(Clk_r), .Q(chosenPacket[26])
         );
  FD4QM1P \Packet_To_Node_reg[26]  ( .D(n34), .CP(Clk_r), .SD(Rst_n), .Q(
        Packet_To_Node[26]) );
  FD1QM1P \chosenPacket_reg[25]  ( .D(n269), .CP(Clk_r), .Q(chosenPacket[25])
         );
  FD2LQM1P \Packet_To_Node_reg[25]  ( .D(n45), .LD(n58), .CP(Clk_r), .CD(Rst_n), .Q(n1) );
  FD1QM1P \chosenPacket_reg[24]  ( .D(n270), .CP(Clk_r), .Q(chosenPacket[24])
         );
  FD1LQM1P \Packet_To_Link_N_reg[31]  ( .D(chosenPacket[31]), .LD(n39), .CP(
        Clk_r), .Q(Packet_To_Link_N[31]) );
  FD1LQM1P \Packet_To_Link_N_reg[30]  ( .D(chosenPacket[30]), .LD(n39), .CP(
        Clk_r), .Q(Packet_To_Link_N[30]) );
  FD1LQM1P \Packet_To_Link_N_reg[29]  ( .D(chosenPacket[29]), .LD(n39), .CP(
        Clk_r), .Q(Packet_To_Link_N[29]) );
  FD1LQM1P \Packet_To_Link_N_reg[27]  ( .D(chosenPacket[27]), .LD(n39), .CP(
        Clk_r), .Q(Packet_To_Link_N[27]) );
  FD1LQM1P \Packet_To_Link_N_reg[25]  ( .D(chosenPacket[25]), .LD(n39), .CP(
        Clk_r), .Q(Packet_To_Link_N[25]) );
  FD1LQM1P \Packet_To_Link_N_reg[16]  ( .D(N108), .LD(n39), .CP(Clk_r), .Q(
        Packet_To_Link_N[16]) );
  FD1LQM1P \Packet_To_Link_N_reg[17]  ( .D(N109), .LD(n39), .CP(Clk_r), .Q(
        Packet_To_Link_N[17]) );
  FD1LQM1P \Packet_To_Link_N_reg[18]  ( .D(N110), .LD(n39), .CP(Clk_r), .Q(
        Packet_To_Link_N[18]) );
  FD1LQM1P \Packet_To_Link_N_reg[19]  ( .D(N111), .LD(n39), .CP(Clk_r), .Q(
        Packet_To_Link_N[19]) );
  FD1LQM1P \Packet_To_Link_N_reg[20]  ( .D(N112), .LD(n39), .CP(Clk_r), .Q(
        Packet_To_Link_N[20]) );
  FD1LQM1P \Packet_To_Link_N_reg[21]  ( .D(N113), .LD(n39), .CP(Clk_r), .Q(
        Packet_To_Link_N[21]) );
  FD1LQM1P \Packet_To_Link_N_reg[22]  ( .D(N114), .LD(n39), .CP(Clk_r), .Q(
        Packet_To_Link_N[22]) );
  FD1LQM1P \Packet_To_Link_N_reg[23]  ( .D(N115), .LD(n39), .CP(Clk_r), .Q(
        Packet_To_Link_N[23]) );
  FD1LQM1P \Packet_To_Link_N_reg[26]  ( .D(chosenPacket[26]), .LD(n39), .CP(
        Clk_r), .Q(Packet_To_Link_N[26]) );
  FD1LQM1P \Packet_To_Link_N_reg[28]  ( .D(chosenPacket[28]), .LD(n39), .CP(
        Clk_r), .Q(Packet_To_Link_N[28]) );
  FD1LQM1P \Packet_To_Link_S_reg[31]  ( .D(chosenPacket[31]), .LD(n40), .CP(
        Clk_r), .Q(Packet_To_Link_S[31]) );
  FD1LQM1P \Packet_To_Link_S_reg[30]  ( .D(chosenPacket[30]), .LD(n40), .CP(
        Clk_r), .Q(Packet_To_Link_S[30]) );
  FD1LQM1P \Packet_To_Link_S_reg[29]  ( .D(chosenPacket[29]), .LD(n40), .CP(
        Clk_r), .Q(Packet_To_Link_S[29]) );
  FD1LQM1P \Packet_To_Link_S_reg[27]  ( .D(chosenPacket[27]), .LD(n40), .CP(
        Clk_r), .Q(Packet_To_Link_S[27]) );
  FD1LQM1P \Packet_To_Link_S_reg[25]  ( .D(chosenPacket[25]), .LD(n40), .CP(
        Clk_r), .Q(Packet_To_Link_S[25]) );
  FD1LQM1P \Packet_To_Link_S_reg[16]  ( .D(N108), .LD(n40), .CP(Clk_r), .Q(
        Packet_To_Link_S[16]) );
  FD1LQM1P \Packet_To_Link_S_reg[17]  ( .D(N109), .LD(n40), .CP(Clk_r), .Q(
        Packet_To_Link_S[17]) );
  FD1LQM1P \Packet_To_Link_S_reg[18]  ( .D(N110), .LD(n40), .CP(Clk_r), .Q(
        Packet_To_Link_S[18]) );
  FD1LQM1P \Packet_To_Link_S_reg[19]  ( .D(N111), .LD(n40), .CP(Clk_r), .Q(
        Packet_To_Link_S[19]) );
  FD1LQM1P \Packet_To_Link_S_reg[20]  ( .D(N112), .LD(n40), .CP(Clk_r), .Q(
        Packet_To_Link_S[20]) );
  FD1LQM1P \Packet_To_Link_S_reg[21]  ( .D(N113), .LD(n40), .CP(Clk_r), .Q(
        Packet_To_Link_S[21]) );
  FD1LQM1P \Packet_To_Link_S_reg[22]  ( .D(N114), .LD(n40), .CP(Clk_r), .Q(
        Packet_To_Link_S[22]) );
  FD1LQM1P \Packet_To_Link_S_reg[23]  ( .D(N115), .LD(n40), .CP(Clk_r), .Q(
        Packet_To_Link_S[23]) );
  FD1LQM1P \Packet_To_Link_S_reg[26]  ( .D(chosenPacket[26]), .LD(n40), .CP(
        Clk_r), .Q(Packet_To_Link_S[26]) );
  FD1LQM1P \Packet_To_Link_S_reg[28]  ( .D(chosenPacket[28]), .LD(n40), .CP(
        Clk_r), .Q(Packet_To_Link_S[28]) );
  FD1LQM1P \Packet_To_Link_W_reg[31]  ( .D(chosenPacket[31]), .LD(n61), .CP(
        Clk_r), .Q(Packet_To_Link_W[31]) );
  FD1LQM1P \Packet_To_Link_W_reg[30]  ( .D(chosenPacket[30]), .LD(n61), .CP(
        Clk_r), .Q(Packet_To_Link_W[30]) );
  FD1LQM1P \Packet_To_Link_W_reg[29]  ( .D(chosenPacket[29]), .LD(n61), .CP(
        Clk_r), .Q(Packet_To_Link_W[29]) );
  FD1LQM1P \Packet_To_Link_W_reg[27]  ( .D(chosenPacket[27]), .LD(n61), .CP(
        Clk_r), .Q(Packet_To_Link_W[27]) );
  FD1LQM1P \Packet_To_Link_W_reg[25]  ( .D(chosenPacket[25]), .LD(n61), .CP(
        Clk_r), .Q(Packet_To_Link_W[25]) );
  FD1LQM1P \Packet_To_Link_W_reg[16]  ( .D(N108), .LD(n61), .CP(Clk_r), .Q(
        Packet_To_Link_W[16]) );
  FD1LQM1P \Packet_To_Link_W_reg[17]  ( .D(N109), .LD(n61), .CP(Clk_r), .Q(
        Packet_To_Link_W[17]) );
  FD1LQM1P \Packet_To_Link_W_reg[18]  ( .D(N110), .LD(n61), .CP(Clk_r), .Q(
        Packet_To_Link_W[18]) );
  FD1LQM1P \Packet_To_Link_W_reg[19]  ( .D(N111), .LD(n61), .CP(Clk_r), .Q(
        Packet_To_Link_W[19]) );
  FD1LQM1P \Packet_To_Link_W_reg[20]  ( .D(N112), .LD(n38), .CP(Clk_r), .Q(
        Packet_To_Link_W[20]) );
  FD1LQM1P \Packet_To_Link_W_reg[21]  ( .D(N113), .LD(n61), .CP(Clk_r), .Q(
        Packet_To_Link_W[21]) );
  FD1LQM1P \Packet_To_Link_W_reg[22]  ( .D(N114), .LD(n61), .CP(Clk_r), .Q(
        Packet_To_Link_W[22]) );
  FD1LQM1P \Packet_To_Link_W_reg[23]  ( .D(N115), .LD(n61), .CP(Clk_r), .Q(
        Packet_To_Link_W[23]) );
  FD1LQM1P \Packet_To_Link_W_reg[26]  ( .D(chosenPacket[26]), .LD(n61), .CP(
        Clk_r), .Q(Packet_To_Link_W[26]) );
  FD1LQM1P \Packet_To_Link_W_reg[28]  ( .D(chosenPacket[28]), .LD(n61), .CP(
        Clk_r), .Q(Packet_To_Link_W[28]) );
  FD1LQM1P \Packet_To_Link_E_reg[31]  ( .D(chosenPacket[31]), .LD(n62), .CP(
        Clk_r), .Q(Packet_To_Link_E[31]) );
  FD1LQM1P \Packet_To_Link_E_reg[30]  ( .D(chosenPacket[30]), .LD(n62), .CP(
        Clk_r), .Q(Packet_To_Link_E[30]) );
  FD1LQM1P \Packet_To_Link_E_reg[29]  ( .D(chosenPacket[29]), .LD(n62), .CP(
        Clk_r), .Q(Packet_To_Link_E[29]) );
  FD1LQM1P \Packet_To_Link_E_reg[27]  ( .D(chosenPacket[27]), .LD(n62), .CP(
        Clk_r), .Q(Packet_To_Link_E[27]) );
  FD1LQM1P \Packet_To_Link_E_reg[25]  ( .D(chosenPacket[25]), .LD(n62), .CP(
        Clk_r), .Q(Packet_To_Link_E[25]) );
  FD1LQM1P \Packet_To_Link_E_reg[16]  ( .D(N108), .LD(n62), .CP(Clk_r), .Q(
        Packet_To_Link_E[16]) );
  FD1LQM1P \Packet_To_Link_E_reg[17]  ( .D(N109), .LD(n62), .CP(Clk_r), .Q(
        Packet_To_Link_E[17]) );
  FD1LQM1P \Packet_To_Link_E_reg[18]  ( .D(N110), .LD(n62), .CP(Clk_r), .Q(
        Packet_To_Link_E[18]) );
  FD1LQM1P \Packet_To_Link_E_reg[19]  ( .D(N111), .LD(n62), .CP(Clk_r), .Q(
        Packet_To_Link_E[19]) );
  FD1LQM1P \Packet_To_Link_E_reg[20]  ( .D(N112), .LD(n62), .CP(Clk_r), .Q(
        Packet_To_Link_E[20]) );
  FD1LQM1P \Packet_To_Link_E_reg[21]  ( .D(N113), .LD(n37), .CP(Clk_r), .Q(
        Packet_To_Link_E[21]) );
  FD1LQM1P \Packet_To_Link_E_reg[22]  ( .D(N114), .LD(n62), .CP(Clk_r), .Q(
        Packet_To_Link_E[22]) );
  FD1LQM1P \Packet_To_Link_E_reg[23]  ( .D(N115), .LD(n62), .CP(Clk_r), .Q(
        Packet_To_Link_E[23]) );
  FD1LQM1P \Packet_To_Link_E_reg[26]  ( .D(chosenPacket[26]), .LD(n62), .CP(
        Clk_r), .Q(Packet_To_Link_E[26]) );
  FD1LQM1P \Packet_To_Link_E_reg[28]  ( .D(chosenPacket[28]), .LD(n62), .CP(
        Clk_r), .Q(Packet_To_Link_E[28]) );
  FD1LQM1P \Packet_To_Link_E_reg[24]  ( .D(chosenPacket[24]), .LD(n62), .CP(
        Clk_r), .Q(Packet_To_Link_E[24]) );
  FD4QM1P \Packet_To_Node_reg[24]  ( .D(n33), .CP(Clk_r), .SD(Rst_n), .Q(
        Packet_To_Node[24]) );
  FD1LQM1P \Packet_To_Link_W_reg[24]  ( .D(chosenPacket[24]), .LD(n61), .CP(
        Clk_r), .Q(Packet_To_Link_W[24]) );
  FD1LQM1P \Packet_To_Link_N_reg[24]  ( .D(chosenPacket[24]), .LD(n39), .CP(
        Clk_r), .Q(Packet_To_Link_N[24]) );
  FD1LQM1P \Packet_To_Link_S_reg[24]  ( .D(chosenPacket[24]), .LD(n40), .CP(
        Clk_r), .Q(Packet_To_Link_S[24]) );
  FD1QM1P \chosenPacket_reg[15]  ( .D(n271), .CP(Clk_r), .Q(chosenPacket[15])
         );
  FD1LQM1P \Packet_To_Link_E_reg[15]  ( .D(chosenPacket[15]), .LD(n62), .CP(
        Clk_r), .Q(Packet_To_Link_E[15]) );
  FD4QM1P \Packet_To_Node_reg[15]  ( .D(n24), .CP(Clk_r), .SD(Rst_n), .Q(
        Packet_To_Node[15]) );
  FD1LQM1P \Packet_To_Link_W_reg[15]  ( .D(chosenPacket[15]), .LD(n61), .CP(
        Clk_r), .Q(Packet_To_Link_W[15]) );
  FD1LQM1P \Packet_To_Link_N_reg[15]  ( .D(chosenPacket[15]), .LD(n39), .CP(
        Clk_r), .Q(Packet_To_Link_N[15]) );
  FD1LQM1P \Packet_To_Link_S_reg[15]  ( .D(chosenPacket[15]), .LD(n40), .CP(
        Clk_r), .Q(Packet_To_Link_S[15]) );
  FD1QM1P \chosenPacket_reg[14]  ( .D(n272), .CP(Clk_r), .Q(chosenPacket[14])
         );
  FD1LQM1P \Packet_To_Link_E_reg[14]  ( .D(chosenPacket[14]), .LD(n62), .CP(
        Clk_r), .Q(Packet_To_Link_E[14]) );
  FD4QM1P \Packet_To_Node_reg[14]  ( .D(n23), .CP(Clk_r), .SD(Rst_n), .Q(
        Packet_To_Node[14]) );
  FD1LQM1P \Packet_To_Link_W_reg[14]  ( .D(chosenPacket[14]), .LD(n61), .CP(
        Clk_r), .Q(Packet_To_Link_W[14]) );
  FD1LQM1P \Packet_To_Link_N_reg[14]  ( .D(chosenPacket[14]), .LD(n39), .CP(
        Clk_r), .Q(Packet_To_Link_N[14]) );
  FD1LQM1P \Packet_To_Link_S_reg[14]  ( .D(chosenPacket[14]), .LD(n40), .CP(
        Clk_r), .Q(Packet_To_Link_S[14]) );
  FD1QM1P \chosenPacket_reg[13]  ( .D(n273), .CP(Clk_r), .Q(chosenPacket[13])
         );
  FD1LQM1P \Packet_To_Link_E_reg[13]  ( .D(chosenPacket[13]), .LD(n62), .CP(
        Clk_r), .Q(Packet_To_Link_E[13]) );
  FD4QM1P \Packet_To_Node_reg[13]  ( .D(n22), .CP(Clk_r), .SD(Rst_n), .Q(
        Packet_To_Node[13]) );
  FD1LQM1P \Packet_To_Link_W_reg[13]  ( .D(chosenPacket[13]), .LD(n61), .CP(
        Clk_r), .Q(Packet_To_Link_W[13]) );
  FD1LQM1P \Packet_To_Link_N_reg[13]  ( .D(chosenPacket[13]), .LD(n39), .CP(
        Clk_r), .Q(Packet_To_Link_N[13]) );
  FD1LQM1P \Packet_To_Link_S_reg[13]  ( .D(chosenPacket[13]), .LD(n40), .CP(
        Clk_r), .Q(Packet_To_Link_S[13]) );
  FD1QM1P \chosenPacket_reg[12]  ( .D(n274), .CP(Clk_r), .Q(chosenPacket[12])
         );
  FD1LQM1P \Packet_To_Link_E_reg[12]  ( .D(chosenPacket[12]), .LD(n62), .CP(
        Clk_r), .Q(Packet_To_Link_E[12]) );
  FD4QM1P \Packet_To_Node_reg[12]  ( .D(n21), .CP(Clk_r), .SD(Rst_n), .Q(
        Packet_To_Node[12]) );
  FD1LQM1P \Packet_To_Link_W_reg[12]  ( .D(chosenPacket[12]), .LD(n61), .CP(
        Clk_r), .Q(Packet_To_Link_W[12]) );
  FD1LQM1P \Packet_To_Link_N_reg[12]  ( .D(chosenPacket[12]), .LD(n39), .CP(
        Clk_r), .Q(Packet_To_Link_N[12]) );
  FD1LQM1P \Packet_To_Link_S_reg[12]  ( .D(chosenPacket[12]), .LD(n40), .CP(
        Clk_r), .Q(Packet_To_Link_S[12]) );
  FD1QM1P \chosenPacket_reg[11]  ( .D(n275), .CP(Clk_r), .Q(chosenPacket[11])
         );
  FD1LQM1P \Packet_To_Link_E_reg[11]  ( .D(chosenPacket[11]), .LD(n62), .CP(
        Clk_r), .Q(Packet_To_Link_E[11]) );
  FD4QM1P \Packet_To_Node_reg[11]  ( .D(n20), .CP(Clk_r), .SD(Rst_n), .Q(
        Packet_To_Node[11]) );
  FD1LQM1P \Packet_To_Link_W_reg[11]  ( .D(chosenPacket[11]), .LD(n61), .CP(
        Clk_r), .Q(Packet_To_Link_W[11]) );
  FD1LQM1P \Packet_To_Link_N_reg[11]  ( .D(chosenPacket[11]), .LD(n39), .CP(
        Clk_r), .Q(Packet_To_Link_N[11]) );
  FD1LQM1P \Packet_To_Link_S_reg[11]  ( .D(chosenPacket[11]), .LD(n40), .CP(
        Clk_r), .Q(Packet_To_Link_S[11]) );
  FD1QM1P \chosenPacket_reg[10]  ( .D(n276), .CP(Clk_r), .Q(chosenPacket[10])
         );
  FD1LQM1P \Packet_To_Link_E_reg[10]  ( .D(chosenPacket[10]), .LD(n62), .CP(
        Clk_r), .Q(Packet_To_Link_E[10]) );
  FD4QM1P \Packet_To_Node_reg[10]  ( .D(n19), .CP(Clk_r), .SD(Rst_n), .Q(
        Packet_To_Node[10]) );
  FD1LQM1P \Packet_To_Link_W_reg[10]  ( .D(chosenPacket[10]), .LD(n38), .CP(
        Clk_r), .Q(Packet_To_Link_W[10]) );
  FD1LQM1P \Packet_To_Link_N_reg[10]  ( .D(chosenPacket[10]), .LD(n39), .CP(
        Clk_r), .Q(Packet_To_Link_N[10]) );
  FD1LQM1P \Packet_To_Link_S_reg[10]  ( .D(chosenPacket[10]), .LD(n40), .CP(
        Clk_r), .Q(Packet_To_Link_S[10]) );
  FD1QM1P \chosenPacket_reg[9]  ( .D(n277), .CP(Clk_r), .Q(chosenPacket[9]) );
  FD1LQM1P \Packet_To_Link_E_reg[9]  ( .D(chosenPacket[9]), .LD(n37), .CP(
        Clk_r), .Q(Packet_To_Link_E[9]) );
  FD4QM1P \Packet_To_Node_reg[9]  ( .D(n18), .CP(Clk_r), .SD(Rst_n), .Q(
        Packet_To_Node[9]) );
  FD1LQM1P \Packet_To_Link_W_reg[9]  ( .D(chosenPacket[9]), .LD(n38), .CP(
        Clk_r), .Q(Packet_To_Link_W[9]) );
  FD1LQM1P \Packet_To_Link_N_reg[9]  ( .D(chosenPacket[9]), .LD(n39), .CP(
        Clk_r), .Q(Packet_To_Link_N[9]) );
  FD1LQM1P \Packet_To_Link_S_reg[9]  ( .D(chosenPacket[9]), .LD(n40), .CP(
        Clk_r), .Q(Packet_To_Link_S[9]) );
  FD1QM1P \chosenPacket_reg[8]  ( .D(n278), .CP(Clk_r), .Q(chosenPacket[8]) );
  FD1LQM1P \Packet_To_Link_E_reg[8]  ( .D(chosenPacket[8]), .LD(n37), .CP(
        Clk_r), .Q(Packet_To_Link_E[8]) );
  FD4QM1P \Packet_To_Node_reg[8]  ( .D(n17), .CP(Clk_r), .SD(Rst_n), .Q(
        Packet_To_Node[8]) );
  FD1LQM1P \Packet_To_Link_W_reg[8]  ( .D(chosenPacket[8]), .LD(n38), .CP(
        Clk_r), .Q(Packet_To_Link_W[8]) );
  FD1LQM1P \Packet_To_Link_N_reg[8]  ( .D(chosenPacket[8]), .LD(n39), .CP(
        Clk_r), .Q(Packet_To_Link_N[8]) );
  FD1LQM1P \Packet_To_Link_S_reg[8]  ( .D(chosenPacket[8]), .LD(n40), .CP(
        Clk_r), .Q(Packet_To_Link_S[8]) );
  FD1QM1P \chosenPacket_reg[7]  ( .D(n279), .CP(Clk_r), .Q(chosenPacket[7]) );
  FD1LQM1P \Packet_To_Link_E_reg[7]  ( .D(chosenPacket[7]), .LD(n37), .CP(
        Clk_r), .Q(Packet_To_Link_E[7]) );
  FD4QM1P \Packet_To_Node_reg[7]  ( .D(n16), .CP(Clk_r), .SD(Rst_n), .Q(
        Packet_To_Node[7]) );
  FD1LQM1P \Packet_To_Link_W_reg[7]  ( .D(chosenPacket[7]), .LD(n38), .CP(
        Clk_r), .Q(Packet_To_Link_W[7]) );
  FD1LQM1P \Packet_To_Link_N_reg[7]  ( .D(chosenPacket[7]), .LD(n39), .CP(
        Clk_r), .Q(Packet_To_Link_N[7]) );
  FD1LQM1P \Packet_To_Link_S_reg[7]  ( .D(chosenPacket[7]), .LD(n40), .CP(
        Clk_r), .Q(Packet_To_Link_S[7]) );
  FD1QM1P \chosenPacket_reg[6]  ( .D(n280), .CP(Clk_r), .Q(chosenPacket[6]) );
  FD1LQM1P \Packet_To_Link_E_reg[6]  ( .D(chosenPacket[6]), .LD(n37), .CP(
        Clk_r), .Q(Packet_To_Link_E[6]) );
  FD4QM1P \Packet_To_Node_reg[6]  ( .D(n15), .CP(Clk_r), .SD(Rst_n), .Q(
        Packet_To_Node[6]) );
  FD1LQM1P \Packet_To_Link_W_reg[6]  ( .D(chosenPacket[6]), .LD(n38), .CP(
        Clk_r), .Q(Packet_To_Link_W[6]) );
  FD1LQM1P \Packet_To_Link_N_reg[6]  ( .D(chosenPacket[6]), .LD(n39), .CP(
        Clk_r), .Q(Packet_To_Link_N[6]) );
  FD1LQM1P \Packet_To_Link_S_reg[6]  ( .D(chosenPacket[6]), .LD(n40), .CP(
        Clk_r), .Q(Packet_To_Link_S[6]) );
  FD1QM1P \chosenPacket_reg[5]  ( .D(n281), .CP(Clk_r), .Q(chosenPacket[5]) );
  FD1LQM1P \Packet_To_Link_E_reg[5]  ( .D(chosenPacket[5]), .LD(n37), .CP(
        Clk_r), .Q(Packet_To_Link_E[5]) );
  FD4QM1P \Packet_To_Node_reg[5]  ( .D(n14), .CP(Clk_r), .SD(Rst_n), .Q(
        Packet_To_Node[5]) );
  FD1LQM1P \Packet_To_Link_W_reg[5]  ( .D(chosenPacket[5]), .LD(n38), .CP(
        Clk_r), .Q(Packet_To_Link_W[5]) );
  FD1LQM1P \Packet_To_Link_N_reg[5]  ( .D(chosenPacket[5]), .LD(n39), .CP(
        Clk_r), .Q(Packet_To_Link_N[5]) );
  FD1LQM1P \Packet_To_Link_S_reg[5]  ( .D(chosenPacket[5]), .LD(n40), .CP(
        Clk_r), .Q(Packet_To_Link_S[5]) );
  FD1QM1P \chosenPacket_reg[4]  ( .D(n282), .CP(Clk_r), .Q(chosenPacket[4]) );
  FD1LQM1P \Packet_To_Link_E_reg[4]  ( .D(chosenPacket[4]), .LD(n37), .CP(
        Clk_r), .Q(Packet_To_Link_E[4]) );
  FD4QM1P \Packet_To_Node_reg[4]  ( .D(n13), .CP(Clk_r), .SD(Rst_n), .Q(
        Packet_To_Node[4]) );
  FD1LQM1P \Packet_To_Link_W_reg[4]  ( .D(chosenPacket[4]), .LD(n61), .CP(
        Clk_r), .Q(Packet_To_Link_W[4]) );
  FD1LQM1P \Packet_To_Link_N_reg[4]  ( .D(chosenPacket[4]), .LD(n39), .CP(
        Clk_r), .Q(Packet_To_Link_N[4]) );
  FD1LQM1P \Packet_To_Link_S_reg[4]  ( .D(chosenPacket[4]), .LD(n40), .CP(
        Clk_r), .Q(Packet_To_Link_S[4]) );
  FD1QM1P \chosenPacket_reg[3]  ( .D(n283), .CP(Clk_r), .Q(chosenPacket[3]) );
  FD1LQM1P \Packet_To_Link_E_reg[3]  ( .D(chosenPacket[3]), .LD(n62), .CP(
        Clk_r), .Q(Packet_To_Link_E[3]) );
  FD4QM1P \Packet_To_Node_reg[3]  ( .D(n12), .CP(Clk_r), .SD(Rst_n), .Q(
        Packet_To_Node[3]) );
  FD1LQM1P \Packet_To_Link_W_reg[3]  ( .D(chosenPacket[3]), .LD(n61), .CP(
        Clk_r), .Q(Packet_To_Link_W[3]) );
  FD1LQM1P \Packet_To_Link_N_reg[3]  ( .D(chosenPacket[3]), .LD(n39), .CP(
        Clk_r), .Q(Packet_To_Link_N[3]) );
  FD1LQM1P \Packet_To_Link_S_reg[3]  ( .D(chosenPacket[3]), .LD(n40), .CP(
        Clk_r), .Q(Packet_To_Link_S[3]) );
  FD1QM1P \chosenPacket_reg[2]  ( .D(n284), .CP(Clk_r), .Q(chosenPacket[2]) );
  FD1LQM1P \Packet_To_Link_E_reg[2]  ( .D(chosenPacket[2]), .LD(n62), .CP(
        Clk_r), .Q(Packet_To_Link_E[2]) );
  FD4QM1P \Packet_To_Node_reg[2]  ( .D(n11), .CP(Clk_r), .SD(Rst_n), .Q(
        Packet_To_Node[2]) );
  FD1LQM1P \Packet_To_Link_W_reg[2]  ( .D(chosenPacket[2]), .LD(n61), .CP(
        Clk_r), .Q(Packet_To_Link_W[2]) );
  FD1LQM1P \Packet_To_Link_N_reg[2]  ( .D(chosenPacket[2]), .LD(n39), .CP(
        Clk_r), .Q(Packet_To_Link_N[2]) );
  FD1LQM1P \Packet_To_Link_S_reg[2]  ( .D(chosenPacket[2]), .LD(n40), .CP(
        Clk_r), .Q(Packet_To_Link_S[2]) );
  FD1QM1P \chosenPacket_reg[1]  ( .D(n285), .CP(Clk_r), .Q(chosenPacket[1]) );
  FD1LQM1P \Packet_To_Link_E_reg[1]  ( .D(chosenPacket[1]), .LD(n62), .CP(
        Clk_r), .Q(Packet_To_Link_E[1]) );
  FD4QM1P \Packet_To_Node_reg[1]  ( .D(n10), .CP(Clk_r), .SD(Rst_n), .Q(
        Packet_To_Node[1]) );
  FD1LQM1P \Packet_To_Link_W_reg[1]  ( .D(chosenPacket[1]), .LD(n61), .CP(
        Clk_r), .Q(Packet_To_Link_W[1]) );
  FD1LQM1P \Packet_To_Link_N_reg[1]  ( .D(chosenPacket[1]), .LD(n39), .CP(
        Clk_r), .Q(Packet_To_Link_N[1]) );
  FD1LQM1P \Packet_To_Link_S_reg[1]  ( .D(chosenPacket[1]), .LD(n40), .CP(
        Clk_r), .Q(Packet_To_Link_S[1]) );
  FD1QM1P \chosenPacket_reg[0]  ( .D(n286), .CP(Clk_r), .Q(chosenPacket[0]) );
  FD1LQM1P \Packet_To_Link_E_reg[0]  ( .D(chosenPacket[0]), .LD(n62), .CP(
        Clk_r), .Q(Packet_To_Link_E[0]) );
  FD4QM1P \Packet_To_Node_reg[0]  ( .D(n9), .CP(Clk_r), .SD(Rst_n), .Q(
        Packet_To_Node[0]) );
  FD1LQM1P \Packet_To_Link_W_reg[0]  ( .D(chosenPacket[0]), .LD(n61), .CP(
        Clk_r), .Q(Packet_To_Link_W[0]) );
  FD1LQM1P \Packet_To_Link_N_reg[0]  ( .D(chosenPacket[0]), .LD(n39), .CP(
        Clk_r), .Q(Packet_To_Link_N[0]) );
  FD1LQM1P \Packet_To_Link_S_reg[0]  ( .D(chosenPacket[0]), .LD(n40), .CP(
        Clk_r), .Q(Packet_To_Link_S[0]) );
  FD1QM1P \chosenPacket_reg[23]  ( .D(n262), .CP(Clk_r), .Q(chosenPacket[23])
         );
  FD1QM1P \chosenPacket_reg[16]  ( .D(n260), .CP(Clk_r), .Q(chosenPacket[16])
         );
  FD1QM1P \chosenPacket_reg[17]  ( .D(n259), .CP(Clk_r), .Q(chosenPacket[17])
         );
  FD1QM1P \chosenPacket_reg[18]  ( .D(n258), .CP(Clk_r), .Q(chosenPacket[18])
         );
  FD1QM1P \chosenPacket_reg[19]  ( .D(n257), .CP(Clk_r), .Q(chosenPacket[19])
         );
  FD1QM1P \chosenPacket_reg[20]  ( .D(n256), .CP(Clk_r), .Q(chosenPacket[20])
         );
  FD1QM1P \chosenPacket_reg[21]  ( .D(n255), .CP(Clk_r), .Q(chosenPacket[21])
         );
  FD1QM1P \chosenPacket_reg[22]  ( .D(n254), .CP(Clk_r), .Q(chosenPacket[22])
         );
  FD4QM1P \RxQueue_Read_reg[1]  ( .D(n218), .CP(Clk_r), .SD(Rst_n), .Q(n50) );
  FD4QM1P \nextStage_reg[0]  ( .D(n7), .CP(Clk_r), .SD(Rst_n), .Q(n8) );
  FD2QM1P \TxQueue_Write_reg[2]  ( .D(n252), .CP(Clk_r), .CD(Rst_n), .Q(
        TxQueue_Write_S) );
  FD2QM1P To_Node_Write_reg ( .D(n261), .CP(Clk_r), .CD(Rst_n), .Q(
        To_Node_Write) );
  FD2QM1P \TxQueue_Write_reg[0]  ( .D(n250), .CP(Clk_r), .CD(Rst_n), .Q(
        TxQueue_Write_E) );
  FD2QM1P \TxQueue_Write_reg[1]  ( .D(n251), .CP(Clk_r), .CD(Rst_n), .Q(
        TxQueue_Write_W) );
  FD2QM1P \RxQueue_Read_reg[2]  ( .D(n247), .CP(Clk_r), .CD(Rst_n), .Q(
        RxQueue_Read_S) );
  FD2QM1P \RxQueue_Read_reg[0]  ( .D(n249), .CP(Clk_r), .CD(Rst_n), .Q(
        RxQueue_Read_E) );
  FD2QM1P \RxQueue_Read_reg[3]  ( .D(n246), .CP(Clk_r), .CD(Rst_n), .Q(
        RxQueue_Read_N) );
  FD2QM1P \RxQueue_Read_reg[4]  ( .D(n245), .CP(Clk_r), .CD(Rst_n), .Q(
        Node_Read) );
  FD2LQM1P \Packet_To_Node_reg[22]  ( .D(n48), .LD(n107), .CP(Clk_r), .CD(
        Rst_n), .Q(n49) );
  FD2QM1P \TxQueue_Write_reg[3]  ( .D(n253), .CP(Clk_r), .CD(Rst_n), .Q(
        TxQueue_Write_N) );
  BUFM1P U3 ( .A(n181), .Z(n53) );
  BUFM1P U4 ( .A(n182), .Z(n54) );
  AOI211M1P U5 ( .A(n43), .B(Router_Address[5]), .C(Router_Address[4]), .D(
        n228), .Z(n31) );
  N1M1P U6 ( .A(n214), .Z(n36) );
  OAI22CDNM1P U7 ( .A(n31), .B(n36), .C(Router_Address[6]), .D(n42), .Z(n46)
         );
  MAJN3M1P U8 ( .A(n41), .B(Router_Address[7]), .C(n46), .Z(n47) );
  ND3CNM1P U9 ( .C(TxQueue_Full_E), .A(Link_Config[0]), .B(n47), .Z(n294) );
  N1M1P U10 ( .A(n49), .Z(Packet_To_Node[22]) );
  N1M1P U11 ( .A(N114), .Z(n48) );
  AND2M4P U12 ( .A(n222), .B(n225), .Z(n40) );
  AND2M4P U13 ( .A(n225), .B(n223), .Z(n39) );
  MUX41HM1P U14 ( .D0(Link_Config[0]), .D1(Link_Config[2]), .D2(Link_Config[1]), .D3(Link_Config[3]), .A(N44), .B(N43), .Z(N48) );
  BUFM1P U15 ( .A(n184), .Z(n56) );
  BUFM1P U16 ( .A(n183), .Z(n55) );
  N1M2P U17 ( .A(n107), .Z(n60) );
  BUFM2P U18 ( .A(n147), .Z(n51) );
  N1M4P U19 ( .A(n50), .Z(RxQueue_Read_W) );
  N1M1P U20 ( .A(n60), .Z(n59) );
  N1M1P U21 ( .A(n60), .Z(n58) );
  BUFM1P U22 ( .A(n148), .Z(n52) );
  NR2M1P U23 ( .A(n219), .B(n51), .Z(n183) );
  NR2BNM1P U24 ( .B(n217), .A(n51), .Z(n182) );
  NR2M1P U25 ( .A(n220), .B(n51), .Z(n181) );
  NR2M1P U26 ( .A(n6), .B(n51), .Z(n184) );
  NR2M1P U27 ( .A(n215), .B(n152), .Z(n297) );
  NR2M1P U28 ( .A(n295), .B(n227), .Z(n38) );
  NR2M1P U29 ( .A(n294), .B(n227), .Z(n37) );
  N1M1P U30 ( .A(chosenPacket[31]), .Z(n41) );
  NR2M1P U31 ( .A(n57), .B(n51), .Z(n148) );
  MUX21LM1P U32 ( .A(chosenPacket[23]), .B(n71), .S(n70), .Z(N115) );
  MUX21LM1P U33 ( .A(chosenPacket[22]), .B(n63), .S(n69), .Z(N114) );
  ND2M1P U34 ( .A(n297), .B(Rst_n), .Z(n147) );
  AND2M1P U35 ( .A(n215), .B(Rst_n), .Z(n225) );
  N1M1P U36 ( .A(n8), .Z(n215) );
  NR2M1P U37 ( .A(dataLocation[0]), .B(n72), .Z(N43) );
  NR2BNM1P U38 ( .B(n299), .A(To_Node_Full), .Z(n107) );
  BUFM2P U39 ( .A(n38), .Z(n61) );
  BUFM2P U40 ( .A(n37), .Z(n62) );
  N1M1P U41 ( .A(n6), .Z(n72) );
  N1M1P U42 ( .A(chosenPacket[22]), .Z(n63) );
  N1M1P U43 ( .A(chosenPacket[20]), .Z(n65) );
  AND3M1P U44 ( .A(chosenPacket[16]), .B(chosenPacket[17]), .C(
        chosenPacket[18]), .Z(n68) );
  ND2M1P U45 ( .A(n68), .B(chosenPacket[19]), .Z(n66) );
  NR2M1P U46 ( .A(n65), .B(n66), .Z(n64) );
  ND2M1P U47 ( .A(n64), .B(chosenPacket[21]), .Z(n69) );
  OR2M1P U48 ( .A(n64), .B(chosenPacket[21]), .Z(n188) );
  ND2M1P U49 ( .A(n69), .B(n188), .Z(n232) );
  N1M1P U50 ( .A(n232), .Z(N113) );
  AOI21M1P U51 ( .A(n66), .B(n65), .C(n64), .Z(N112) );
  OAI21M1P U52 ( .A(n68), .B(chosenPacket[19]), .C(n66), .Z(n234) );
  N1M1P U53 ( .A(n234), .Z(N111) );
  AOI21M1P U54 ( .A(chosenPacket[17]), .B(chosenPacket[16]), .C(
        chosenPacket[18]), .Z(n67) );
  NR2M1P U55 ( .A(n68), .B(n67), .Z(N110) );
  OAI22CDNM1P U56 ( .A(chosenPacket[17]), .B(chosenPacket[16]), .C(
        chosenPacket[16]), .D(chosenPacket[17]), .Z(n236) );
  N1M1P U57 ( .A(n236), .Z(N109) );
  N1M1P U58 ( .A(chosenPacket[16]), .Z(N108) );
  N1M1P U59 ( .A(chosenPacket[23]), .Z(n71) );
  ND2BNM1P U60 ( .B(n69), .A(chosenPacket[22]), .Z(n70) );
  N1M1P U61 ( .A(chosenPacket[25]), .Z(n45) );
  N1M1P U62 ( .A(chosenPacket[27]), .Z(n44) );
  N1M1P U63 ( .A(chosenPacket[29]), .Z(n43) );
  N1M1P U64 ( .A(chosenPacket[30]), .Z(n42) );
  ND3M1P U65 ( .A(dataLocation[0]), .B(n6), .C(dataLocation[1]), .Z(n57) );
  ND2M1P U66 ( .A(N43), .B(dataLocation[1]), .Z(n220) );
  NR3CNM1P U67 ( .C(dataLocation[0]), .A(dataLocation[1]), .B(n72), .Z(n73) );
  N1M1P U68 ( .A(n73), .Z(n219) );
  ND2M1P U69 ( .A(n220), .B(n219), .Z(N44) );
  AOI22DNM1P U70 ( .A(RxQueue_Empty_E), .B(n72), .D(N48), .C(n57), .Z(n76) );
  AOI22DNM1P U71 ( .A(n73), .B(RxQueue_Empty_S), .D(n57), .C(Node_Queue_Empty), 
        .Z(n75) );
  NR2BNM1P U72 ( .B(N43), .A(dataLocation[1]), .Z(n217) );
  AOI22DNM1P U73 ( .A(n217), .B(RxQueue_Empty_W), .D(n220), .C(RxQueue_Empty_N), .Z(n74) );
  ND3M1P U74 ( .A(n76), .B(n75), .C(n74), .Z(n152) );
  AOI22M1P U75 ( .A(Packet_From_Link_E[0]), .B(n56), .C(chosenPacket[0]), .D(
        n51), .Z(n79) );
  AOI22M1P U76 ( .A(n181), .B(Packet_From_Link_N[0]), .C(n183), .D(
        Packet_From_Link_S[0]), .Z(n78) );
  AOI22M1P U77 ( .A(n54), .B(Packet_From_Link_W[0]), .C(n148), .D(
        Packet_From_Node[0]), .Z(n77) );
  ND3M1P U78 ( .A(n79), .B(n78), .C(n77), .Z(n286) );
  AOI22M1P U79 ( .A(Packet_From_Link_E[1]), .B(n56), .C(chosenPacket[1]), .D(
        n51), .Z(n82) );
  AOI22M1P U80 ( .A(n181), .B(Packet_From_Link_N[1]), .C(n183), .D(
        Packet_From_Link_S[1]), .Z(n81) );
  AOI22M1P U81 ( .A(n54), .B(Packet_From_Link_W[1]), .C(n148), .D(
        Packet_From_Node[1]), .Z(n80) );
  ND3M1P U82 ( .A(n82), .B(n81), .C(n80), .Z(n285) );
  AOI22M1P U83 ( .A(Packet_From_Link_E[2]), .B(n184), .C(chosenPacket[2]), .D(
        n51), .Z(n85) );
  AOI22M1P U84 ( .A(n181), .B(Packet_From_Link_N[2]), .C(n183), .D(
        Packet_From_Link_S[2]), .Z(n84) );
  AOI22M1P U85 ( .A(n54), .B(Packet_From_Link_W[2]), .C(n148), .D(
        Packet_From_Node[2]), .Z(n83) );
  ND3M1P U86 ( .A(n85), .B(n84), .C(n83), .Z(n284) );
  AOI22M1P U87 ( .A(Packet_From_Link_E[3]), .B(n56), .C(chosenPacket[3]), .D(
        n51), .Z(n88) );
  AOI22M1P U88 ( .A(n181), .B(Packet_From_Link_N[3]), .C(n183), .D(
        Packet_From_Link_S[3]), .Z(n87) );
  AOI22M1P U89 ( .A(n54), .B(Packet_From_Link_W[3]), .C(n148), .D(
        Packet_From_Node[3]), .Z(n86) );
  ND3M1P U90 ( .A(n88), .B(n87), .C(n86), .Z(n283) );
  AOI22M1P U91 ( .A(Packet_From_Link_E[4]), .B(n56), .C(chosenPacket[4]), .D(
        n51), .Z(n91) );
  AOI22M1P U92 ( .A(n181), .B(Packet_From_Link_N[4]), .C(n183), .D(
        Packet_From_Link_S[4]), .Z(n90) );
  AOI22M1P U93 ( .A(n54), .B(Packet_From_Link_W[4]), .C(n148), .D(
        Packet_From_Node[4]), .Z(n89) );
  ND3M1P U94 ( .A(n91), .B(n90), .C(n89), .Z(n282) );
  AOI22M1P U95 ( .A(Packet_From_Link_E[5]), .B(n56), .C(chosenPacket[5]), .D(
        n51), .Z(n94) );
  AOI22M1P U96 ( .A(n181), .B(Packet_From_Link_N[5]), .C(n183), .D(
        Packet_From_Link_S[5]), .Z(n93) );
  AOI22M1P U97 ( .A(n182), .B(Packet_From_Link_W[5]), .C(n148), .D(
        Packet_From_Node[5]), .Z(n92) );
  ND3M1P U98 ( .A(n94), .B(n93), .C(n92), .Z(n281) );
  AOI22M1P U99 ( .A(Packet_From_Link_E[6]), .B(n56), .C(chosenPacket[6]), .D(
        n51), .Z(n97) );
  AOI22M1P U100 ( .A(n181), .B(Packet_From_Link_N[6]), .C(n183), .D(
        Packet_From_Link_S[6]), .Z(n96) );
  AOI22M1P U101 ( .A(n182), .B(Packet_From_Link_W[6]), .C(n148), .D(
        Packet_From_Node[6]), .Z(n95) );
  ND3M1P U102 ( .A(n97), .B(n96), .C(n95), .Z(n280) );
  AOI22M1P U103 ( .A(Packet_From_Link_E[7]), .B(n56), .C(chosenPacket[7]), .D(
        n51), .Z(n100) );
  AOI22M1P U104 ( .A(n181), .B(Packet_From_Link_N[7]), .C(n183), .D(
        Packet_From_Link_S[7]), .Z(n99) );
  AOI22M1P U105 ( .A(n182), .B(Packet_From_Link_W[7]), .C(n148), .D(
        Packet_From_Node[7]), .Z(n98) );
  ND3M1P U106 ( .A(n100), .B(n99), .C(n98), .Z(n279) );
  AOI22M1P U107 ( .A(Packet_From_Link_E[8]), .B(n184), .C(chosenPacket[8]), 
        .D(n51), .Z(n103) );
  AOI22M1P U108 ( .A(n53), .B(Packet_From_Link_N[8]), .C(n55), .D(
        Packet_From_Link_S[8]), .Z(n102) );
  AOI22M1P U109 ( .A(n54), .B(Packet_From_Link_W[8]), .C(n52), .D(
        Packet_From_Node[8]), .Z(n101) );
  ND3M1P U110 ( .A(n103), .B(n102), .C(n101), .Z(n278) );
  AOI22M1P U111 ( .A(Packet_From_Link_E[9]), .B(n56), .C(chosenPacket[9]), .D(
        n51), .Z(n106) );
  AOI22M1P U112 ( .A(n53), .B(Packet_From_Link_N[9]), .C(n183), .D(
        Packet_From_Link_S[9]), .Z(n105) );
  AOI22M1P U113 ( .A(n54), .B(Packet_From_Link_W[9]), .C(n52), .D(
        Packet_From_Node[9]), .Z(n104) );
  ND3M1P U114 ( .A(n106), .B(n105), .C(n104), .Z(n277) );
  AOI22M1P U115 ( .A(Packet_From_Link_E[10]), .B(n184), .C(chosenPacket[10]), 
        .D(n51), .Z(n110) );
  AOI22M1P U116 ( .A(n53), .B(Packet_From_Link_N[10]), .C(n55), .D(
        Packet_From_Link_S[10]), .Z(n109) );
  AOI22M1P U117 ( .A(n182), .B(Packet_From_Link_W[10]), .C(n52), .D(
        Packet_From_Node[10]), .Z(n108) );
  ND3M1P U118 ( .A(n110), .B(n109), .C(n108), .Z(n276) );
  AOI22M1P U119 ( .A(Packet_From_Link_E[11]), .B(n56), .C(chosenPacket[11]), 
        .D(n51), .Z(n113) );
  AOI22M1P U120 ( .A(n53), .B(Packet_From_Link_N[11]), .C(n55), .D(
        Packet_From_Link_S[11]), .Z(n112) );
  AOI22M1P U121 ( .A(n54), .B(Packet_From_Link_W[11]), .C(n52), .D(
        Packet_From_Node[11]), .Z(n111) );
  ND3M1P U122 ( .A(n113), .B(n112), .C(n111), .Z(n275) );
  AOI22M1P U123 ( .A(Packet_From_Link_E[12]), .B(n184), .C(chosenPacket[12]), 
        .D(n51), .Z(n116) );
  AOI22M1P U124 ( .A(n53), .B(Packet_From_Link_N[12]), .C(n55), .D(
        Packet_From_Link_S[12]), .Z(n115) );
  AOI22M1P U125 ( .A(n182), .B(Packet_From_Link_W[12]), .C(n52), .D(
        Packet_From_Node[12]), .Z(n114) );
  ND3M1P U126 ( .A(n116), .B(n115), .C(n114), .Z(n274) );
  AOI22M1P U127 ( .A(Packet_From_Link_E[13]), .B(n184), .C(chosenPacket[13]), 
        .D(n51), .Z(n119) );
  AOI22M1P U128 ( .A(n53), .B(Packet_From_Link_N[13]), .C(n55), .D(
        Packet_From_Link_S[13]), .Z(n118) );
  AOI22M1P U129 ( .A(n54), .B(Packet_From_Link_W[13]), .C(n52), .D(
        Packet_From_Node[13]), .Z(n117) );
  ND3M1P U130 ( .A(n119), .B(n118), .C(n117), .Z(n273) );
  AOI22M1P U131 ( .A(Packet_From_Link_E[14]), .B(n184), .C(chosenPacket[14]), 
        .D(n51), .Z(n122) );
  AOI22M1P U132 ( .A(n53), .B(Packet_From_Link_N[14]), .C(n55), .D(
        Packet_From_Link_S[14]), .Z(n121) );
  AOI22M1P U133 ( .A(n182), .B(Packet_From_Link_W[14]), .C(n52), .D(
        Packet_From_Node[14]), .Z(n120) );
  ND3M1P U134 ( .A(n122), .B(n121), .C(n120), .Z(n272) );
  AOI22M1P U135 ( .A(Packet_From_Link_E[15]), .B(n184), .C(chosenPacket[15]), 
        .D(n51), .Z(n125) );
  AOI22M1P U136 ( .A(n53), .B(Packet_From_Link_N[15]), .C(n55), .D(
        Packet_From_Link_S[15]), .Z(n124) );
  AOI22M1P U137 ( .A(n54), .B(Packet_From_Link_W[15]), .C(n52), .D(
        Packet_From_Node[15]), .Z(n123) );
  ND3M1P U138 ( .A(n125), .B(n124), .C(n123), .Z(n271) );
  AOI22M1P U139 ( .A(chosenPacket[24]), .B(n51), .C(n184), .D(
        Packet_From_Link_E[24]), .Z(n128) );
  AOI22M1P U140 ( .A(n181), .B(Packet_From_Link_N[24]), .C(n183), .D(
        Packet_From_Link_S[24]), .Z(n127) );
  AOI22M1P U141 ( .A(n54), .B(Packet_From_Link_W[24]), .C(n52), .D(
        Packet_From_Node_24), .Z(n126) );
  ND3M1P U142 ( .A(n128), .B(n127), .C(n126), .Z(n270) );
  AOI22M1P U143 ( .A(chosenPacket[25]), .B(n51), .C(n184), .D(
        Packet_From_Link_E[25]), .Z(n131) );
  AOI22M1P U144 ( .A(n181), .B(Packet_From_Link_N[25]), .C(n183), .D(
        Packet_From_Link_S[25]), .Z(n130) );
  AOI22M1P U145 ( .A(n54), .B(Packet_From_Link_W[25]), .C(n52), .D(
        Packet_From_Node_25), .Z(n129) );
  ND3M1P U146 ( .A(n131), .B(n130), .C(n129), .Z(n269) );
  AOI22M1P U147 ( .A(chosenPacket[26]), .B(n51), .C(n184), .D(
        Packet_From_Link_E[26]), .Z(n134) );
  AOI22M1P U148 ( .A(n181), .B(Packet_From_Link_N[26]), .C(n183), .D(
        Packet_From_Link_S[26]), .Z(n133) );
  AOI22M1P U149 ( .A(n54), .B(Packet_From_Link_W[26]), .C(n52), .D(
        Packet_From_Node_26), .Z(n132) );
  ND3M1P U150 ( .A(n134), .B(n133), .C(n132), .Z(n268) );
  AOI22M1P U151 ( .A(chosenPacket[27]), .B(n51), .C(n56), .D(
        Packet_From_Link_E[27]), .Z(n137) );
  AOI22M1P U152 ( .A(n53), .B(Packet_From_Link_N[27]), .C(n55), .D(
        Packet_From_Link_S[27]), .Z(n136) );
  AOI22M1P U153 ( .A(n182), .B(Packet_From_Link_W[27]), .C(n52), .D(
        Packet_From_Node_27), .Z(n135) );
  ND3M1P U154 ( .A(n137), .B(n136), .C(n135), .Z(n267) );
  AOI22M1P U155 ( .A(chosenPacket[28]), .B(n51), .C(n184), .D(
        Packet_From_Link_E[28]), .Z(n140) );
  AOI22M1P U156 ( .A(n53), .B(Packet_From_Link_N[28]), .C(n55), .D(
        Packet_From_Link_S[28]), .Z(n139) );
  AOI22M1P U157 ( .A(n54), .B(Packet_From_Link_W[28]), .C(n148), .D(
        Packet_From_Node_28), .Z(n138) );
  ND3M1P U158 ( .A(n140), .B(n139), .C(n138), .Z(n266) );
  AOI22M1P U159 ( .A(chosenPacket[29]), .B(n147), .C(n184), .D(
        Packet_From_Link_E[29]), .Z(n143) );
  AOI22M1P U160 ( .A(n53), .B(Packet_From_Link_N[29]), .C(n55), .D(
        Packet_From_Link_S[29]), .Z(n142) );
  AOI22M1P U161 ( .A(n54), .B(Packet_From_Link_W[29]), .C(n52), .D(
        Packet_From_Node_29), .Z(n141) );
  ND3M1P U162 ( .A(n143), .B(n142), .C(n141), .Z(n265) );
  AOI22M1P U163 ( .A(chosenPacket[30]), .B(n147), .C(n56), .D(
        Packet_From_Link_E[30]), .Z(n146) );
  AOI22M1P U164 ( .A(n53), .B(Packet_From_Link_N[30]), .C(n55), .D(
        Packet_From_Link_S[30]), .Z(n145) );
  AOI22M1P U165 ( .A(n54), .B(Packet_From_Link_W[30]), .C(n148), .D(
        Packet_From_Node_30), .Z(n144) );
  ND3M1P U166 ( .A(n146), .B(n145), .C(n144), .Z(n264) );
  AOI22M1P U167 ( .A(chosenPacket[31]), .B(n51), .C(n56), .D(
        Packet_From_Link_E[31]), .Z(n151) );
  AOI22M1P U168 ( .A(n53), .B(Packet_From_Link_N[31]), .C(n55), .D(
        Packet_From_Link_S[31]), .Z(n150) );
  AOI22M1P U169 ( .A(n54), .B(Packet_From_Link_W[31]), .C(n52), .D(
        Packet_From_Node_31), .Z(n149) );
  ND3M1P U170 ( .A(n151), .B(n150), .C(n149), .Z(n263) );
  AO21CNM1P U171 ( .A(n8), .B(n152), .C(Rst_n), .Z(n180) );
  AOI22M1P U172 ( .A(chosenPacket[23]), .B(n180), .C(N115), .D(n225), .Z(n155)
         );
  AOI22M1P U173 ( .A(n54), .B(Packet_From_Link_W[23]), .C(n53), .D(
        Packet_From_Link_N[23]), .Z(n154) );
  AOI22M1P U174 ( .A(n56), .B(Packet_From_Link_E[23]), .C(n55), .D(
        Packet_From_Link_S[23]), .Z(n153) );
  ND3M1P U175 ( .A(n155), .B(n154), .C(n153), .Z(n262) );
  N1M1P U176 ( .A(chosenPacket[24]), .Z(n230) );
  N1M1P U177 ( .A(chosenPacket[28]), .Z(n228) );
  ND2M1P U178 ( .A(Router_Address[3]), .B(n44), .Z(n204) );
  ND2M1P U179 ( .A(Router_Address[4]), .B(n228), .Z(n208) );
  OAI211M1P U180 ( .A(Router_Address[4]), .B(n228), .C(n204), .D(n208), .Z(
        n159) );
  NR2M1P U181 ( .A(Router_Address[5]), .B(n43), .Z(n207) );
  NR2M1P U182 ( .A(Router_Address[6]), .B(n42), .Z(n210) );
  NR2M1P U183 ( .A(n207), .B(n210), .Z(n214) );
  AOI22M1P U184 ( .A(Router_Address[5]), .B(n43), .C(Router_Address[6]), .D(
        n42), .Z(n206) );
  NR2M1P U185 ( .A(Router_Address[3]), .B(n44), .Z(n156) );
  NR2M1P U186 ( .A(Router_Address[0]), .B(n230), .Z(n193) );
  AOI211M1P U187 ( .A(Router_Address[1]), .B(n45), .C(n156), .D(n193), .Z(n157) );
  N1M1P U188 ( .A(chosenPacket[26]), .Z(n229) );
  ND2M1P U189 ( .A(Router_Address[2]), .B(n229), .Z(n192) );
  ND4M1P U190 ( .A(n214), .B(n206), .C(n157), .D(n192), .Z(n158) );
  AOI211M1P U191 ( .A(Router_Address[0]), .B(n230), .C(n159), .D(n158), .Z(
        n161) );
  OAI22M1P U192 ( .A(Router_Address[2]), .B(n229), .C(Router_Address[1]), .D(
        n45), .Z(n198) );
  AOI21M1P U193 ( .A(Router_Address[7]), .B(n41), .C(n198), .Z(n160) );
  OAI211M1P U194 ( .A(Router_Address[7]), .B(n41), .C(n161), .D(n160), .Z(n189) );
  NR2M1P U195 ( .A(n8), .B(n189), .Z(n299) );
  AO21CNM1P U196 ( .A(To_Node_Write), .B(n215), .C(n60), .Z(n261) );
  AOI22M1P U197 ( .A(chosenPacket[16]), .B(n180), .C(n225), .D(N108), .Z(n164)
         );
  AOI22M1P U198 ( .A(n56), .B(Packet_From_Link_E[16]), .C(n53), .D(
        Packet_From_Link_N[16]), .Z(n163) );
  AOI22M1P U199 ( .A(n54), .B(Packet_From_Link_W[16]), .C(n55), .D(
        Packet_From_Link_S[16]), .Z(n162) );
  ND3M1P U200 ( .A(n164), .B(n163), .C(n162), .Z(n260) );
  AOI22M1P U201 ( .A(chosenPacket[17]), .B(n180), .C(n225), .D(N109), .Z(n167)
         );
  AOI22M1P U202 ( .A(n54), .B(Packet_From_Link_W[17]), .C(n53), .D(
        Packet_From_Link_N[17]), .Z(n166) );
  AOI22M1P U203 ( .A(n56), .B(Packet_From_Link_E[17]), .C(n55), .D(
        Packet_From_Link_S[17]), .Z(n165) );
  ND3M1P U204 ( .A(n167), .B(n166), .C(n165), .Z(n259) );
  AOI22M1P U205 ( .A(chosenPacket[18]), .B(n180), .C(n225), .D(N110), .Z(n170)
         );
  AOI22M1P U206 ( .A(n54), .B(Packet_From_Link_W[18]), .C(n53), .D(
        Packet_From_Link_N[18]), .Z(n169) );
  AOI22M1P U207 ( .A(n56), .B(Packet_From_Link_E[18]), .C(n55), .D(
        Packet_From_Link_S[18]), .Z(n168) );
  ND3M1P U208 ( .A(n170), .B(n169), .C(n168), .Z(n258) );
  AOI22M1P U209 ( .A(chosenPacket[19]), .B(n180), .C(N111), .D(n225), .Z(n173)
         );
  AOI22M1P U210 ( .A(n54), .B(Packet_From_Link_W[19]), .C(n53), .D(
        Packet_From_Link_N[19]), .Z(n172) );
  AOI22M1P U211 ( .A(n56), .B(Packet_From_Link_E[19]), .C(n55), .D(
        Packet_From_Link_S[19]), .Z(n171) );
  ND3M1P U212 ( .A(n173), .B(n172), .C(n171), .Z(n257) );
  AOI22M1P U213 ( .A(chosenPacket[20]), .B(n180), .C(N112), .D(n225), .Z(n176)
         );
  AOI22M1P U214 ( .A(n54), .B(Packet_From_Link_W[20]), .C(n53), .D(
        Packet_From_Link_N[20]), .Z(n175) );
  AOI22M1P U215 ( .A(n56), .B(Packet_From_Link_E[20]), .C(n55), .D(
        Packet_From_Link_S[20]), .Z(n174) );
  ND3M1P U216 ( .A(n176), .B(n175), .C(n174), .Z(n256) );
  AOI22M1P U217 ( .A(chosenPacket[21]), .B(n180), .C(n225), .D(N113), .Z(n179)
         );
  AOI22M1P U218 ( .A(n182), .B(Packet_From_Link_W[21]), .C(n53), .D(
        Packet_From_Link_N[21]), .Z(n178) );
  AOI22M1P U219 ( .A(n56), .B(Packet_From_Link_E[21]), .C(n55), .D(
        Packet_From_Link_S[21]), .Z(n177) );
  ND3M1P U220 ( .A(n179), .B(n178), .C(n177), .Z(n255) );
  AOI22M1P U221 ( .A(chosenPacket[22]), .B(n180), .C(N114), .D(n225), .Z(n187)
         );
  AOI22M1P U222 ( .A(n182), .B(Packet_From_Link_W[22]), .C(n53), .D(
        Packet_From_Link_N[22]), .Z(n186) );
  AOI22M1P U223 ( .A(n56), .B(Packet_From_Link_E[22]), .C(n55), .D(
        Packet_From_Link_S[22]), .Z(n185) );
  ND3M1P U224 ( .A(n187), .B(n186), .C(n185), .Z(n254) );
  ND4M1P U225 ( .A(chosenPacket[17]), .B(chosenPacket[18]), .C(
        chosenPacket[19]), .D(N108), .Z(n191) );
  ND4M1P U226 ( .A(N115), .B(N114), .C(N112), .D(n188), .Z(n190) );
  OA21M1P U227 ( .A(n191), .B(n190), .C(n189), .Z(n197) );
  N1M1P U228 ( .A(n192), .Z(n202) );
  ND2M1P U229 ( .A(Router_Address[1]), .B(n45), .Z(n200) );
  AOI21M1P U230 ( .A(n193), .B(n200), .C(n198), .Z(n194) );
  OAI22M1P U231 ( .A(n202), .B(n194), .C(Router_Address[3]), .D(n44), .Z(n195)
         );
  ND4DNM1P U232 ( .D(TxQueue_Full_N), .A(Link_Config[3]), .B(n195), .C(n204), 
        .Z(n196) );
  NR2BNM1P U233 ( .B(n197), .A(n196), .Z(n223) );
  OA21M1P U234 ( .A(n223), .B(TxQueue_Write_N), .C(n215), .Z(n253) );
  ND2M1P U235 ( .A(n197), .B(n196), .Z(n226) );
  ND2M1P U236 ( .A(Router_Address[0]), .B(n230), .Z(n199) );
  AOI21M1P U237 ( .A(n200), .B(n199), .C(n198), .Z(n201) );
  OAI22M1P U238 ( .A(n202), .B(n201), .C(Router_Address[3]), .D(n44), .Z(n203)
         );
  AOI21M1P U239 ( .A(n204), .B(n203), .C(TxQueue_Full_S), .Z(n205) );
  ND2M1P U240 ( .A(Link_Config[2]), .B(n205), .Z(n224) );
  NR2M1P U241 ( .A(n226), .B(n224), .Z(n222) );
  OA21M1P U242 ( .A(n222), .B(TxQueue_Write_S), .C(n215), .Z(n252) );
  N1M1P U243 ( .A(Router_Address[7]), .Z(n212) );
  OAI21M1P U244 ( .A(n208), .B(n207), .C(n206), .Z(n209) );
  ND2BNM1P U245 ( .B(n210), .A(n209), .Z(n211) );
  MAJN3M1P U246 ( .A(chosenPacket[31]), .B(n212), .C(n211), .Z(n213) );
  ND3CNM1P U247 ( .C(TxQueue_Full_W), .A(Link_Config[1]), .B(n213), .Z(n295)
         );
  NR3CNM1P U248 ( .C(n224), .A(n226), .B(n8), .Z(n296) );
  N1M1P U249 ( .A(n296), .Z(n216) );
  OAI22CDNM1P U250 ( .A(n295), .B(n216), .C(n215), .D(TxQueue_Write_W), .Z(
        n251) );
  OAI22CDNM1P U251 ( .A(n294), .B(n216), .C(n215), .D(TxQueue_Write_E), .Z(
        n250) );
  N1M1P U252 ( .A(n297), .Z(n221) );
  OAI22CDNM1P U253 ( .A(n6), .B(n221), .C(n8), .D(RxQueue_Read_E), .Z(n249) );
  AOI22M1P U254 ( .A(n8), .B(RxQueue_Read_W), .C(n217), .D(n297), .Z(n218) );
  OAI22CDNM1P U255 ( .A(n219), .B(n221), .C(n8), .D(RxQueue_Read_S), .Z(n247)
         );
  OAI22CDNM1P U256 ( .A(n220), .B(n221), .C(n8), .D(RxQueue_Read_N), .Z(n246)
         );
  OAI22CDNM1P U257 ( .A(n57), .B(n221), .C(n8), .D(Node_Read), .Z(n245) );
  ND3CNM1P U258 ( .C(n226), .A(n225), .B(n224), .Z(n227) );
  AOI22DNM1P U259 ( .A(n58), .B(n228), .D(Packet_To_Node[28]), .C(n60), .Z(n35) );
  AOI22DNM1P U260 ( .A(n58), .B(n229), .D(Packet_To_Node[26]), .C(n60), .Z(n34) );
  AOI22DNM1P U261 ( .A(n58), .B(n230), .D(Packet_To_Node[24]), .C(n60), .Z(n33) );
  OAI22M1P U262 ( .A(n60), .B(N115), .C(Packet_To_Node[23]), .D(n58), .Z(n231)
         );
  N1M1P U263 ( .A(n231), .Z(n32) );
  AOI22DNM1P U264 ( .A(n58), .B(n232), .D(Packet_To_Node[21]), .C(n60), .Z(n30) );
  OAI22M1P U265 ( .A(n60), .B(N112), .C(Packet_To_Node[20]), .D(n59), .Z(n233)
         );
  N1M1P U266 ( .A(n233), .Z(n29) );
  AOI22DNM1P U267 ( .A(n58), .B(n234), .D(Packet_To_Node[19]), .C(n60), .Z(n28) );
  OAI22M1P U268 ( .A(n60), .B(N110), .C(Packet_To_Node[18]), .D(n59), .Z(n235)
         );
  N1M1P U269 ( .A(n235), .Z(n27) );
  AOI22DNM1P U270 ( .A(n58), .B(n236), .D(Packet_To_Node[17]), .C(n60), .Z(n26) );
  AOI22DNM1P U271 ( .A(n58), .B(chosenPacket[16]), .D(Packet_To_Node[16]), .C(
        n60), .Z(n25) );
  OAI22M1P U272 ( .A(n60), .B(chosenPacket[15]), .C(Packet_To_Node[15]), .D(
        n59), .Z(n237) );
  N1M1P U273 ( .A(n237), .Z(n24) );
  OAI22M1P U274 ( .A(n60), .B(chosenPacket[14]), .C(Packet_To_Node[14]), .D(
        n59), .Z(n238) );
  N1M1P U275 ( .A(n238), .Z(n23) );
  OAI22M1P U276 ( .A(n60), .B(chosenPacket[13]), .C(Packet_To_Node[13]), .D(
        n59), .Z(n239) );
  N1M1P U277 ( .A(n239), .Z(n22) );
  OAI22M1P U278 ( .A(n60), .B(chosenPacket[12]), .C(Packet_To_Node[12]), .D(
        n59), .Z(n240) );
  N1M1P U279 ( .A(n240), .Z(n21) );
  OAI22M1P U280 ( .A(n60), .B(chosenPacket[11]), .C(Packet_To_Node[11]), .D(
        n59), .Z(n241) );
  N1M1P U281 ( .A(n241), .Z(n20) );
  OAI22M1P U282 ( .A(n60), .B(chosenPacket[10]), .C(Packet_To_Node[10]), .D(
        n59), .Z(n242) );
  N1M1P U283 ( .A(n242), .Z(n19) );
  OAI22M1P U284 ( .A(n60), .B(chosenPacket[9]), .C(Packet_To_Node[9]), .D(n59), 
        .Z(n243) );
  N1M1P U285 ( .A(n243), .Z(n18) );
  OAI22M1P U286 ( .A(n60), .B(chosenPacket[8]), .C(Packet_To_Node[8]), .D(n59), 
        .Z(n244) );
  N1M1P U287 ( .A(n244), .Z(n17) );
  OAI22M1P U288 ( .A(n60), .B(chosenPacket[7]), .C(Packet_To_Node[7]), .D(n59), 
        .Z(n248) );
  N1M1P U289 ( .A(n248), .Z(n16) );
  OAI22M1P U290 ( .A(n60), .B(chosenPacket[6]), .C(Packet_To_Node[6]), .D(n59), 
        .Z(n287) );
  N1M1P U291 ( .A(n287), .Z(n15) );
  OAI22M1P U292 ( .A(n60), .B(chosenPacket[5]), .C(Packet_To_Node[5]), .D(n59), 
        .Z(n288) );
  N1M1P U293 ( .A(n288), .Z(n14) );
  OAI22M1P U294 ( .A(n60), .B(chosenPacket[4]), .C(Packet_To_Node[4]), .D(n59), 
        .Z(n289) );
  N1M1P U295 ( .A(n289), .Z(n13) );
  OAI22M1P U296 ( .A(n60), .B(chosenPacket[3]), .C(Packet_To_Node[3]), .D(n59), 
        .Z(n290) );
  N1M1P U297 ( .A(n290), .Z(n12) );
  OAI22M1P U298 ( .A(n60), .B(chosenPacket[2]), .C(Packet_To_Node[2]), .D(n59), 
        .Z(n291) );
  N1M1P U299 ( .A(n291), .Z(n11) );
  OAI22M1P U300 ( .A(n60), .B(chosenPacket[1]), .C(Packet_To_Node[1]), .D(n59), 
        .Z(n292) );
  N1M1P U301 ( .A(n292), .Z(n10) );
  OAI22M1P U302 ( .A(n60), .B(chosenPacket[0]), .C(Packet_To_Node[0]), .D(n58), 
        .Z(n293) );
  N1M1P U303 ( .A(n293), .Z(n9) );
  AND3M1P U304 ( .A(n296), .B(n295), .C(n294), .Z(n298) );
  AOI211M1P U305 ( .A(To_Node_Full), .B(n299), .C(n298), .D(n297), .Z(n7) );
  N1M1P U306 ( .A(n5), .Z(Packet_To_Node[31]) );
  N1M1P U307 ( .A(n4), .Z(Packet_To_Node[30]) );
  N1M1P U308 ( .A(n3), .Z(Packet_To_Node[29]) );
  N1M1P U309 ( .A(n2), .Z(Packet_To_Node[27]) );
  N1M1P U310 ( .A(n1), .Z(Packet_To_Node[25]) );
endmodule


module Packet_Queue_1 ( Clk_r, Rst_n, Packet_In, Read_Ack, Write_Ack, 
        Packet_Out, Empty, Full );
  input [31:0] Packet_In;
  output [31:0] Packet_Out;
  input Clk_r, Rst_n, Read_Ack, Write_Ack;
  output Empty, Full;
  wire   \Queue[4][31] , \Queue[4][30] , \Queue[4][29] , \Queue[4][28] ,
         \Queue[4][27] , \Queue[4][26] , \Queue[4][25] , \Queue[4][24] ,
         \Queue[4][23] , \Queue[4][22] , \Queue[4][21] , \Queue[4][20] ,
         \Queue[4][19] , \Queue[4][18] , \Queue[4][17] , \Queue[4][16] ,
         \Queue[4][15] , \Queue[4][14] , \Queue[4][13] , \Queue[4][12] ,
         \Queue[4][11] , \Queue[4][10] , \Queue[4][9] , \Queue[4][8] ,
         \Queue[4][7] , \Queue[4][6] , \Queue[4][5] , \Queue[4][4] ,
         \Queue[4][3] , \Queue[4][2] , \Queue[4][1] , \Queue[4][0] ,
         \Queue[3][31] , \Queue[3][30] , \Queue[3][29] , \Queue[3][28] ,
         \Queue[3][27] , \Queue[3][26] , \Queue[3][25] , \Queue[3][24] ,
         \Queue[3][23] , \Queue[3][22] , \Queue[3][21] , \Queue[3][20] ,
         \Queue[3][19] , \Queue[3][18] , \Queue[3][17] , \Queue[3][16] ,
         \Queue[3][15] , \Queue[3][14] , \Queue[3][13] , \Queue[3][12] ,
         \Queue[3][11] , \Queue[3][10] , \Queue[3][9] , \Queue[3][8] ,
         \Queue[3][7] , \Queue[3][6] , \Queue[3][5] , \Queue[3][4] ,
         \Queue[3][3] , \Queue[3][2] , \Queue[3][1] , \Queue[3][0] ,
         \Queue[2][31] , \Queue[2][30] , \Queue[2][29] , \Queue[2][28] ,
         \Queue[2][27] , \Queue[2][26] , \Queue[2][25] , \Queue[2][24] ,
         \Queue[2][23] , \Queue[2][22] , \Queue[2][21] , \Queue[2][20] ,
         \Queue[2][19] , \Queue[2][18] , \Queue[2][17] , \Queue[2][16] ,
         \Queue[2][15] , \Queue[2][14] , \Queue[2][13] , \Queue[2][12] ,
         \Queue[2][11] , \Queue[2][10] , \Queue[2][9] , \Queue[2][8] ,
         \Queue[2][7] , \Queue[2][6] , \Queue[2][5] , \Queue[2][4] ,
         \Queue[2][3] , \Queue[2][2] , \Queue[2][1] , \Queue[2][0] ,
         \Queue[1][31] , \Queue[1][30] , \Queue[1][29] , \Queue[1][28] ,
         \Queue[1][27] , \Queue[1][26] , \Queue[1][25] , \Queue[1][24] ,
         \Queue[1][23] , \Queue[1][22] , \Queue[1][21] , \Queue[1][20] ,
         \Queue[1][19] , \Queue[1][18] , \Queue[1][17] , \Queue[1][16] ,
         \Queue[1][15] , \Queue[1][14] , \Queue[1][13] , \Queue[1][12] ,
         \Queue[1][11] , \Queue[1][10] , \Queue[1][9] , \Queue[1][8] ,
         \Queue[1][7] , \Queue[1][6] , \Queue[1][5] , \Queue[1][4] ,
         \Queue[1][3] , \Queue[1][2] , \Queue[1][1] , \Queue[1][0] , n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534;
  wire   [2:0] Count;

  FDN2QM1P \Count_reg[0]  ( .D(n207), .CPN(Clk_r), .CD(Rst_n), .Q(Count[0]) );
  FDN2QM1P \Count_reg[1]  ( .D(n208), .CPN(Clk_r), .CD(Rst_n), .Q(Count[1]) );
  FDN2QM1P \Count_reg[2]  ( .D(n371), .CPN(Clk_r), .CD(Rst_n), .Q(Count[2]) );
  FDN1QM1P \Queue_reg[4][30]  ( .D(n403), .CPN(Clk_r), .Q(\Queue[4][30] ) );
  FDN1QM1P \Queue_reg[3][30]  ( .D(n531), .CPN(Clk_r), .Q(\Queue[3][30] ) );
  FDN1QM1P \Queue_reg[2][30]  ( .D(n499), .CPN(Clk_r), .Q(\Queue[2][30] ) );
  FDN1QM1P \Queue_reg[4][29]  ( .D(n402), .CPN(Clk_r), .Q(\Queue[4][29] ) );
  FDN1QM1P \Queue_reg[3][29]  ( .D(n530), .CPN(Clk_r), .Q(\Queue[3][29] ) );
  FDN1QM1P \Queue_reg[2][29]  ( .D(n498), .CPN(Clk_r), .Q(\Queue[2][29] ) );
  FDN1QM1P \Queue_reg[4][28]  ( .D(n401), .CPN(Clk_r), .Q(\Queue[4][28] ) );
  FDN1QM1P \Queue_reg[3][28]  ( .D(n529), .CPN(Clk_r), .Q(\Queue[3][28] ) );
  FDN1QM1P \Queue_reg[2][28]  ( .D(n497), .CPN(Clk_r), .Q(\Queue[2][28] ) );
  FDN1QM1P \Queue_reg[4][27]  ( .D(n400), .CPN(Clk_r), .Q(\Queue[4][27] ) );
  FDN1QM1P \Queue_reg[3][27]  ( .D(n528), .CPN(Clk_r), .Q(\Queue[3][27] ) );
  FDN1QM1P \Queue_reg[2][27]  ( .D(n496), .CPN(Clk_r), .Q(\Queue[2][27] ) );
  FDN1QM1P \Queue_reg[4][26]  ( .D(n399), .CPN(Clk_r), .Q(\Queue[4][26] ) );
  FDN1QM1P \Queue_reg[3][26]  ( .D(n527), .CPN(Clk_r), .Q(\Queue[3][26] ) );
  FDN1QM1P \Queue_reg[2][26]  ( .D(n495), .CPN(Clk_r), .Q(\Queue[2][26] ) );
  FDN1QM1P \Queue_reg[4][25]  ( .D(n398), .CPN(Clk_r), .Q(\Queue[4][25] ) );
  FDN1QM1P \Queue_reg[3][25]  ( .D(n526), .CPN(Clk_r), .Q(\Queue[3][25] ) );
  FDN1QM1P \Queue_reg[2][25]  ( .D(n494), .CPN(Clk_r), .Q(\Queue[2][25] ) );
  FDN1QM1P \Queue_reg[4][24]  ( .D(n397), .CPN(Clk_r), .Q(\Queue[4][24] ) );
  FDN1QM1P \Queue_reg[3][24]  ( .D(n525), .CPN(Clk_r), .Q(\Queue[3][24] ) );
  FDN1QM1P \Queue_reg[2][24]  ( .D(n493), .CPN(Clk_r), .Q(\Queue[2][24] ) );
  FDN1QM1P \Queue_reg[4][23]  ( .D(n396), .CPN(Clk_r), .Q(\Queue[4][23] ) );
  FDN1QM1P \Queue_reg[3][23]  ( .D(n524), .CPN(Clk_r), .Q(\Queue[3][23] ) );
  FDN1QM1P \Queue_reg[2][23]  ( .D(n492), .CPN(Clk_r), .Q(\Queue[2][23] ) );
  FDN1QM1P \Queue_reg[4][22]  ( .D(n395), .CPN(Clk_r), .Q(\Queue[4][22] ) );
  FDN1QM1P \Queue_reg[3][22]  ( .D(n523), .CPN(Clk_r), .Q(\Queue[3][22] ) );
  FDN1QM1P \Queue_reg[2][22]  ( .D(n491), .CPN(Clk_r), .Q(\Queue[2][22] ) );
  FDN1QM1P \Queue_reg[4][21]  ( .D(n394), .CPN(Clk_r), .Q(\Queue[4][21] ) );
  FDN1QM1P \Queue_reg[3][21]  ( .D(n522), .CPN(Clk_r), .Q(\Queue[3][21] ) );
  FDN1QM1P \Queue_reg[2][21]  ( .D(n490), .CPN(Clk_r), .Q(\Queue[2][21] ) );
  FDN1QM1P \Queue_reg[4][20]  ( .D(n393), .CPN(Clk_r), .Q(\Queue[4][20] ) );
  FDN1QM1P \Queue_reg[3][20]  ( .D(n521), .CPN(Clk_r), .Q(\Queue[3][20] ) );
  FDN1QM1P \Queue_reg[2][20]  ( .D(n489), .CPN(Clk_r), .Q(\Queue[2][20] ) );
  FDN1QM1P \Queue_reg[4][19]  ( .D(n392), .CPN(Clk_r), .Q(\Queue[4][19] ) );
  FDN1QM1P \Queue_reg[3][19]  ( .D(n520), .CPN(Clk_r), .Q(\Queue[3][19] ) );
  FDN1QM1P \Queue_reg[2][19]  ( .D(n488), .CPN(Clk_r), .Q(\Queue[2][19] ) );
  FDN1QM1P \Queue_reg[4][18]  ( .D(n391), .CPN(Clk_r), .Q(\Queue[4][18] ) );
  FDN1QM1P \Queue_reg[3][18]  ( .D(n519), .CPN(Clk_r), .Q(\Queue[3][18] ) );
  FDN1QM1P \Queue_reg[2][18]  ( .D(n487), .CPN(Clk_r), .Q(\Queue[2][18] ) );
  FDN1QM1P \Queue_reg[4][17]  ( .D(n390), .CPN(Clk_r), .Q(\Queue[4][17] ) );
  FDN1QM1P \Queue_reg[3][17]  ( .D(n518), .CPN(Clk_r), .Q(\Queue[3][17] ) );
  FDN1QM1P \Queue_reg[2][17]  ( .D(n486), .CPN(Clk_r), .Q(\Queue[2][17] ) );
  FDN1QM1P \Queue_reg[4][16]  ( .D(n389), .CPN(Clk_r), .Q(\Queue[4][16] ) );
  FDN1QM1P \Queue_reg[3][16]  ( .D(n517), .CPN(Clk_r), .Q(\Queue[3][16] ) );
  FDN1QM1P \Queue_reg[2][16]  ( .D(n485), .CPN(Clk_r), .Q(\Queue[2][16] ) );
  FDN1QM1P \Queue_reg[4][15]  ( .D(n388), .CPN(Clk_r), .Q(\Queue[4][15] ) );
  FDN1QM1P \Queue_reg[3][15]  ( .D(n516), .CPN(Clk_r), .Q(\Queue[3][15] ) );
  FDN1QM1P \Queue_reg[2][15]  ( .D(n484), .CPN(Clk_r), .Q(\Queue[2][15] ) );
  FDN1QM1P \Queue_reg[4][14]  ( .D(n387), .CPN(Clk_r), .Q(\Queue[4][14] ) );
  FDN1QM1P \Queue_reg[3][14]  ( .D(n515), .CPN(Clk_r), .Q(\Queue[3][14] ) );
  FDN1QM1P \Queue_reg[2][14]  ( .D(n483), .CPN(Clk_r), .Q(\Queue[2][14] ) );
  FDN1QM1P \Queue_reg[4][13]  ( .D(n386), .CPN(Clk_r), .Q(\Queue[4][13] ) );
  FDN1QM1P \Queue_reg[3][13]  ( .D(n514), .CPN(Clk_r), .Q(\Queue[3][13] ) );
  FDN1QM1P \Queue_reg[2][13]  ( .D(n482), .CPN(Clk_r), .Q(\Queue[2][13] ) );
  FDN1QM1P \Queue_reg[4][12]  ( .D(n385), .CPN(Clk_r), .Q(\Queue[4][12] ) );
  FDN1QM1P \Queue_reg[3][12]  ( .D(n513), .CPN(Clk_r), .Q(\Queue[3][12] ) );
  FDN1QM1P \Queue_reg[2][12]  ( .D(n481), .CPN(Clk_r), .Q(\Queue[2][12] ) );
  FDN1QM1P \Queue_reg[4][11]  ( .D(n384), .CPN(Clk_r), .Q(\Queue[4][11] ) );
  FDN1QM1P \Queue_reg[3][11]  ( .D(n512), .CPN(Clk_r), .Q(\Queue[3][11] ) );
  FDN1QM1P \Queue_reg[2][11]  ( .D(n480), .CPN(Clk_r), .Q(\Queue[2][11] ) );
  FDN1QM1P \Queue_reg[4][10]  ( .D(n383), .CPN(Clk_r), .Q(\Queue[4][10] ) );
  FDN1QM1P \Queue_reg[3][10]  ( .D(n511), .CPN(Clk_r), .Q(\Queue[3][10] ) );
  FDN1QM1P \Queue_reg[2][10]  ( .D(n479), .CPN(Clk_r), .Q(\Queue[2][10] ) );
  FDN1QM1P \Queue_reg[4][9]  ( .D(n382), .CPN(Clk_r), .Q(\Queue[4][9] ) );
  FDN1QM1P \Queue_reg[3][9]  ( .D(n510), .CPN(Clk_r), .Q(\Queue[3][9] ) );
  FDN1QM1P \Queue_reg[2][9]  ( .D(n478), .CPN(Clk_r), .Q(\Queue[2][9] ) );
  FDN1QM1P \Queue_reg[4][8]  ( .D(n381), .CPN(Clk_r), .Q(\Queue[4][8] ) );
  FDN1QM1P \Queue_reg[3][8]  ( .D(n509), .CPN(Clk_r), .Q(\Queue[3][8] ) );
  FDN1QM1P \Queue_reg[2][8]  ( .D(n477), .CPN(Clk_r), .Q(\Queue[2][8] ) );
  FDN1QM1P \Queue_reg[4][7]  ( .D(n380), .CPN(Clk_r), .Q(\Queue[4][7] ) );
  FDN1QM1P \Queue_reg[3][7]  ( .D(n508), .CPN(Clk_r), .Q(\Queue[3][7] ) );
  FDN1QM1P \Queue_reg[2][7]  ( .D(n476), .CPN(Clk_r), .Q(\Queue[2][7] ) );
  FDN1QM1P \Queue_reg[4][6]  ( .D(n379), .CPN(Clk_r), .Q(\Queue[4][6] ) );
  FDN1QM1P \Queue_reg[3][6]  ( .D(n507), .CPN(Clk_r), .Q(\Queue[3][6] ) );
  FDN1QM1P \Queue_reg[2][6]  ( .D(n475), .CPN(Clk_r), .Q(\Queue[2][6] ) );
  FDN1QM1P \Queue_reg[4][5]  ( .D(n378), .CPN(Clk_r), .Q(\Queue[4][5] ) );
  FDN1QM1P \Queue_reg[3][5]  ( .D(n506), .CPN(Clk_r), .Q(\Queue[3][5] ) );
  FDN1QM1P \Queue_reg[2][5]  ( .D(n474), .CPN(Clk_r), .Q(\Queue[2][5] ) );
  FDN1QM1P \Queue_reg[4][4]  ( .D(n377), .CPN(Clk_r), .Q(\Queue[4][4] ) );
  FDN1QM1P \Queue_reg[3][4]  ( .D(n505), .CPN(Clk_r), .Q(\Queue[3][4] ) );
  FDN1QM1P \Queue_reg[2][4]  ( .D(n473), .CPN(Clk_r), .Q(\Queue[2][4] ) );
  FDN1QM1P \Queue_reg[4][3]  ( .D(n376), .CPN(Clk_r), .Q(\Queue[4][3] ) );
  FDN1QM1P \Queue_reg[3][3]  ( .D(n504), .CPN(Clk_r), .Q(\Queue[3][3] ) );
  FDN1QM1P \Queue_reg[2][3]  ( .D(n472), .CPN(Clk_r), .Q(\Queue[2][3] ) );
  FDN1QM1P \Queue_reg[4][2]  ( .D(n375), .CPN(Clk_r), .Q(\Queue[4][2] ) );
  FDN1QM1P \Queue_reg[3][2]  ( .D(n503), .CPN(Clk_r), .Q(\Queue[3][2] ) );
  FDN1QM1P \Queue_reg[2][2]  ( .D(n471), .CPN(Clk_r), .Q(\Queue[2][2] ) );
  FDN1QM1P \Queue_reg[4][1]  ( .D(n374), .CPN(Clk_r), .Q(\Queue[4][1] ) );
  FDN1QM1P \Queue_reg[3][1]  ( .D(n502), .CPN(Clk_r), .Q(\Queue[3][1] ) );
  FDN1QM1P \Queue_reg[2][1]  ( .D(n470), .CPN(Clk_r), .Q(\Queue[2][1] ) );
  FDN1QM1P \Queue_reg[4][0]  ( .D(n373), .CPN(Clk_r), .Q(\Queue[4][0] ) );
  FDN1QM1P \Queue_reg[3][0]  ( .D(n501), .CPN(Clk_r), .Q(\Queue[3][0] ) );
  FDN1QM1P \Queue_reg[2][0]  ( .D(n469), .CPN(Clk_r), .Q(\Queue[2][0] ) );
  FDN1QM1P \Queue_reg[4][31]  ( .D(n372), .CPN(Clk_r), .Q(\Queue[4][31] ) );
  FDN1QM1P \Queue_reg[3][31]  ( .D(n532), .CPN(Clk_r), .Q(\Queue[3][31] ) );
  FDN1QM1P \Queue_reg[2][31]  ( .D(n500), .CPN(Clk_r), .Q(\Queue[2][31] ) );
  FDN2QM1P Full_reg ( .D(n404), .CPN(Clk_r), .CD(Rst_n), .Q(Full) );
  FDN1QM1P \Queue_reg[1][31]  ( .D(n436), .CPN(Clk_r), .Q(\Queue[1][31] ) );
  FDN1QM1P \Queue_reg[0][31]  ( .D(n468), .CPN(Clk_r), .Q(Packet_Out[31]) );
  FDN1QM1P \Queue_reg[1][30]  ( .D(n435), .CPN(Clk_r), .Q(\Queue[1][30] ) );
  FDN1QM1P \Queue_reg[0][30]  ( .D(n467), .CPN(Clk_r), .Q(Packet_Out[30]) );
  FDN1QM1P \Queue_reg[1][29]  ( .D(n434), .CPN(Clk_r), .Q(\Queue[1][29] ) );
  FDN1QM1P \Queue_reg[0][29]  ( .D(n466), .CPN(Clk_r), .Q(Packet_Out[29]) );
  FDN1QM1P \Queue_reg[1][28]  ( .D(n433), .CPN(Clk_r), .Q(\Queue[1][28] ) );
  FDN1QM1P \Queue_reg[0][28]  ( .D(n465), .CPN(Clk_r), .Q(Packet_Out[28]) );
  FDN1QM1P \Queue_reg[1][27]  ( .D(n432), .CPN(Clk_r), .Q(\Queue[1][27] ) );
  FDN1QM1P \Queue_reg[0][27]  ( .D(n464), .CPN(Clk_r), .Q(Packet_Out[27]) );
  FDN1QM1P \Queue_reg[1][26]  ( .D(n431), .CPN(Clk_r), .Q(\Queue[1][26] ) );
  FDN1QM1P \Queue_reg[0][26]  ( .D(n463), .CPN(Clk_r), .Q(Packet_Out[26]) );
  FDN1QM1P \Queue_reg[1][25]  ( .D(n430), .CPN(Clk_r), .Q(\Queue[1][25] ) );
  FDN1QM1P \Queue_reg[0][25]  ( .D(n462), .CPN(Clk_r), .Q(Packet_Out[25]) );
  FDN1QM1P \Queue_reg[1][24]  ( .D(n429), .CPN(Clk_r), .Q(\Queue[1][24] ) );
  FDN1QM1P \Queue_reg[0][24]  ( .D(n461), .CPN(Clk_r), .Q(Packet_Out[24]) );
  FDN1QM1P \Queue_reg[1][23]  ( .D(n428), .CPN(Clk_r), .Q(\Queue[1][23] ) );
  FDN1QM1P \Queue_reg[0][23]  ( .D(n460), .CPN(Clk_r), .Q(Packet_Out[23]) );
  FDN1QM1P \Queue_reg[1][22]  ( .D(n427), .CPN(Clk_r), .Q(\Queue[1][22] ) );
  FDN1QM1P \Queue_reg[0][22]  ( .D(n459), .CPN(Clk_r), .Q(Packet_Out[22]) );
  FDN1QM1P \Queue_reg[1][21]  ( .D(n426), .CPN(Clk_r), .Q(\Queue[1][21] ) );
  FDN1QM1P \Queue_reg[0][21]  ( .D(n458), .CPN(Clk_r), .Q(Packet_Out[21]) );
  FDN1QM1P \Queue_reg[1][20]  ( .D(n425), .CPN(Clk_r), .Q(\Queue[1][20] ) );
  FDN1QM1P \Queue_reg[0][20]  ( .D(n457), .CPN(Clk_r), .Q(Packet_Out[20]) );
  FDN1QM1P \Queue_reg[1][19]  ( .D(n424), .CPN(Clk_r), .Q(\Queue[1][19] ) );
  FDN1QM1P \Queue_reg[0][19]  ( .D(n456), .CPN(Clk_r), .Q(Packet_Out[19]) );
  FDN1QM1P \Queue_reg[1][18]  ( .D(n423), .CPN(Clk_r), .Q(\Queue[1][18] ) );
  FDN1QM1P \Queue_reg[0][18]  ( .D(n455), .CPN(Clk_r), .Q(Packet_Out[18]) );
  FDN1QM1P \Queue_reg[1][17]  ( .D(n422), .CPN(Clk_r), .Q(\Queue[1][17] ) );
  FDN1QM1P \Queue_reg[0][17]  ( .D(n454), .CPN(Clk_r), .Q(Packet_Out[17]) );
  FDN1QM1P \Queue_reg[1][16]  ( .D(n421), .CPN(Clk_r), .Q(\Queue[1][16] ) );
  FDN1QM1P \Queue_reg[0][16]  ( .D(n453), .CPN(Clk_r), .Q(Packet_Out[16]) );
  FDN1QM1P \Queue_reg[1][15]  ( .D(n420), .CPN(Clk_r), .Q(\Queue[1][15] ) );
  FDN1QM1P \Queue_reg[0][15]  ( .D(n452), .CPN(Clk_r), .Q(Packet_Out[15]) );
  FDN1QM1P \Queue_reg[1][14]  ( .D(n419), .CPN(Clk_r), .Q(\Queue[1][14] ) );
  FDN1QM1P \Queue_reg[0][14]  ( .D(n451), .CPN(Clk_r), .Q(Packet_Out[14]) );
  FDN1QM1P \Queue_reg[1][13]  ( .D(n418), .CPN(Clk_r), .Q(\Queue[1][13] ) );
  FDN1QM1P \Queue_reg[0][13]  ( .D(n450), .CPN(Clk_r), .Q(Packet_Out[13]) );
  FDN1QM1P \Queue_reg[1][12]  ( .D(n417), .CPN(Clk_r), .Q(\Queue[1][12] ) );
  FDN1QM1P \Queue_reg[0][12]  ( .D(n449), .CPN(Clk_r), .Q(Packet_Out[12]) );
  FDN1QM1P \Queue_reg[1][11]  ( .D(n416), .CPN(Clk_r), .Q(\Queue[1][11] ) );
  FDN1QM1P \Queue_reg[0][11]  ( .D(n448), .CPN(Clk_r), .Q(Packet_Out[11]) );
  FDN1QM1P \Queue_reg[1][10]  ( .D(n415), .CPN(Clk_r), .Q(\Queue[1][10] ) );
  FDN1QM1P \Queue_reg[0][10]  ( .D(n447), .CPN(Clk_r), .Q(Packet_Out[10]) );
  FDN1QM1P \Queue_reg[1][9]  ( .D(n414), .CPN(Clk_r), .Q(\Queue[1][9] ) );
  FDN1QM1P \Queue_reg[0][9]  ( .D(n446), .CPN(Clk_r), .Q(Packet_Out[9]) );
  FDN1QM1P \Queue_reg[1][8]  ( .D(n413), .CPN(Clk_r), .Q(\Queue[1][8] ) );
  FDN1QM1P \Queue_reg[0][8]  ( .D(n445), .CPN(Clk_r), .Q(Packet_Out[8]) );
  FDN1QM1P \Queue_reg[1][7]  ( .D(n412), .CPN(Clk_r), .Q(\Queue[1][7] ) );
  FDN1QM1P \Queue_reg[0][7]  ( .D(n444), .CPN(Clk_r), .Q(Packet_Out[7]) );
  FDN1QM1P \Queue_reg[1][6]  ( .D(n411), .CPN(Clk_r), .Q(\Queue[1][6] ) );
  FDN1QM1P \Queue_reg[0][6]  ( .D(n443), .CPN(Clk_r), .Q(Packet_Out[6]) );
  FDN1QM1P \Queue_reg[1][5]  ( .D(n410), .CPN(Clk_r), .Q(\Queue[1][5] ) );
  FDN1QM1P \Queue_reg[0][5]  ( .D(n442), .CPN(Clk_r), .Q(Packet_Out[5]) );
  FDN1QM1P \Queue_reg[1][4]  ( .D(n409), .CPN(Clk_r), .Q(\Queue[1][4] ) );
  FDN1QM1P \Queue_reg[0][4]  ( .D(n441), .CPN(Clk_r), .Q(Packet_Out[4]) );
  FDN1QM1P \Queue_reg[1][3]  ( .D(n408), .CPN(Clk_r), .Q(\Queue[1][3] ) );
  FDN1QM1P \Queue_reg[0][3]  ( .D(n440), .CPN(Clk_r), .Q(Packet_Out[3]) );
  FDN1QM1P \Queue_reg[1][2]  ( .D(n407), .CPN(Clk_r), .Q(\Queue[1][2] ) );
  FDN1QM1P \Queue_reg[0][2]  ( .D(n439), .CPN(Clk_r), .Q(Packet_Out[2]) );
  FDN1QM1P \Queue_reg[1][1]  ( .D(n406), .CPN(Clk_r), .Q(\Queue[1][1] ) );
  FDN1QM1P \Queue_reg[0][1]  ( .D(n438), .CPN(Clk_r), .Q(Packet_Out[1]) );
  FDN1QM1P \Queue_reg[1][0]  ( .D(n405), .CPN(Clk_r), .Q(\Queue[1][0] ) );
  FDN1QM1P \Queue_reg[0][0]  ( .D(n437), .CPN(Clk_r), .Q(Packet_Out[0]) );
  FDN2QM1P Empty_reg ( .D(n534), .CPN(Clk_r), .CD(Rst_n), .Q(n533) );
  NR3M1P U3 ( .A(Count[0]), .B(Count[2]), .C(n16), .Z(n94) );
  N1M1P U4 ( .A(Read_Ack), .Z(n131) );
  N1M1P U5 ( .A(n3), .Z(n93) );
  NR3M1P U6 ( .A(n17), .B(Count[2]), .C(Count[1]), .Z(n206) );
  NR3M1P U7 ( .A(Count[2]), .B(n17), .C(n16), .Z(n134) );
  AOI21M3P U8 ( .A(n3), .B(n94), .C(n135), .Z(n51) );
  OAI211M4P U9 ( .A(n94), .B(n131), .C(n3), .D(n18), .Z(n53) );
  OAI211M4P U10 ( .A(n206), .B(n131), .C(n3), .D(n56), .Z(n91) );
  AOI21M3P U11 ( .A(n3), .B(n136), .C(n135), .Z(n199) );
  AOI21M3P U12 ( .A(n3), .B(n134), .C(n135), .Z(n126) );
  NR2FM3P U13 ( .A(n55), .B(n15), .Z(n14) );
  OAI211M4P U14 ( .A(n94), .B(n133), .C(Rst_n), .D(n132), .Z(n127) );
  OAI211M4P U15 ( .A(n134), .B(n133), .C(Rst_n), .D(n132), .Z(n200) );
  OAI211M4P U16 ( .A(n136), .B(n131), .C(n3), .D(n130), .Z(n202) );
  OAI211M4P U17 ( .A(n134), .B(n131), .C(n3), .D(n92), .Z(n129) );
  OAI21M2P U18 ( .A(n3), .B(Read_Ack), .C(n18), .Z(n50) );
  N1M1P U19 ( .A(n136), .Z(n15) );
  NR3M1P U20 ( .A(Count[0]), .B(Count[1]), .C(n13), .Z(n136) );
  N1M1P U21 ( .A(Count[1]), .Z(n16) );
  N1M1P U22 ( .A(Count[2]), .Z(n13) );
  N1M1P U23 ( .A(Count[0]), .Z(n17) );
  N1M3P U24 ( .A(n12), .Z(n133) );
  BUFM3P U25 ( .A(n89), .Z(n6) );
  ND2M2P U26 ( .A(Read_Ack), .B(Rst_n), .Z(n135) );
  ND2M2P U27 ( .A(n12), .B(Rst_n), .Z(n55) );
  NR2FM2P U28 ( .A(Read_Ack), .B(n93), .Z(n12) );
  BUFM10P U29 ( .A(Write_Ack), .Z(n3) );
  N1M1P U30 ( .A(Packet_In[25]), .Z(n188) );
  N1M1P U31 ( .A(Packet_In[31]), .Z(n203) );
  N1M1P U32 ( .A(Packet_In[27]), .Z(n192) );
  N1M1P U33 ( .A(Packet_In[29]), .Z(n196) );
  N1M1P U34 ( .A(Packet_In[30]), .Z(n198) );
  BUFM2P U35 ( .A(n50), .Z(n4) );
  BUFM2P U36 ( .A(n50), .Z(n5) );
  N1M2P U37 ( .A(n56), .Z(n88) );
  NR2M1P U38 ( .A(n131), .B(n3), .Z(n205) );
  NR2M1P U39 ( .A(n12), .B(n205), .Z(n204) );
  AOI22CDNM1P U40 ( .A(n204), .B(n17), .C(n204), .D(n17), .Z(n207) );
  N1M1P U41 ( .A(n205), .Z(n11) );
  AOI22M1P U42 ( .A(Count[0]), .B(n133), .C(n11), .D(n17), .Z(n8) );
  AOI22CDNM1P U43 ( .A(Count[1]), .B(n8), .C(n8), .D(Count[1]), .Z(n208) );
  ND3M1P U44 ( .A(n17), .B(n13), .C(n16), .Z(n54) );
  ND2M1P U45 ( .A(Count[1]), .B(Read_Ack), .Z(n7) );
  OAI211M1P U46 ( .A(Count[1]), .B(n133), .C(n8), .D(n7), .Z(n9) );
  AOI22M1P U47 ( .A(n12), .B(n134), .C(Count[2]), .D(n9), .Z(n10) );
  OAI21M1P U48 ( .A(n54), .B(n11), .C(n10), .Z(n371) );
  AOI22CDNM1P U49 ( .A(n14), .B(n203), .C(\Queue[4][31] ), .D(n14), .Z(n372)
         );
  N1M1P U50 ( .A(Packet_In[0]), .Z(n138) );
  AOI22CDNM1P U51 ( .A(n14), .B(n138), .C(\Queue[4][0] ), .D(n14), .Z(n373) );
  N1M1P U52 ( .A(Packet_In[1]), .Z(n140) );
  AOI22CDNM1P U53 ( .A(n14), .B(n140), .C(\Queue[4][1] ), .D(n14), .Z(n374) );
  N1M1P U54 ( .A(Packet_In[2]), .Z(n142) );
  AOI22CDNM1P U55 ( .A(n14), .B(n142), .C(\Queue[4][2] ), .D(n14), .Z(n375) );
  N1M1P U56 ( .A(Packet_In[3]), .Z(n144) );
  AOI22CDNM1P U57 ( .A(n14), .B(n144), .C(\Queue[4][3] ), .D(n14), .Z(n376) );
  N1M1P U58 ( .A(Packet_In[4]), .Z(n146) );
  AOI22CDNM1P U59 ( .A(n14), .B(n146), .C(\Queue[4][4] ), .D(n14), .Z(n377) );
  N1M1P U60 ( .A(Packet_In[5]), .Z(n148) );
  AOI22CDNM1P U61 ( .A(n14), .B(n148), .C(\Queue[4][5] ), .D(n14), .Z(n378) );
  N1M1P U62 ( .A(Packet_In[6]), .Z(n150) );
  AOI22CDNM1P U63 ( .A(n14), .B(n150), .C(\Queue[4][6] ), .D(n14), .Z(n379) );
  N1M1P U64 ( .A(Packet_In[7]), .Z(n152) );
  AOI22CDNM1P U65 ( .A(n14), .B(n152), .C(\Queue[4][7] ), .D(n14), .Z(n380) );
  N1M1P U66 ( .A(Packet_In[8]), .Z(n154) );
  AOI22CDNM1P U67 ( .A(n14), .B(n154), .C(\Queue[4][8] ), .D(n14), .Z(n381) );
  N1M1P U68 ( .A(Packet_In[9]), .Z(n156) );
  AOI22CDNM1P U69 ( .A(n14), .B(n156), .C(\Queue[4][9] ), .D(n14), .Z(n382) );
  N1M1P U70 ( .A(Packet_In[10]), .Z(n158) );
  AOI22CDNM1P U71 ( .A(n14), .B(n158), .C(\Queue[4][10] ), .D(n14), .Z(n383)
         );
  N1M1P U72 ( .A(Packet_In[11]), .Z(n160) );
  AOI22CDNM1P U73 ( .A(n14), .B(n160), .C(\Queue[4][11] ), .D(n14), .Z(n384)
         );
  N1M1P U74 ( .A(Packet_In[12]), .Z(n162) );
  AOI22CDNM1P U75 ( .A(n14), .B(n162), .C(\Queue[4][12] ), .D(n14), .Z(n385)
         );
  N1M1P U76 ( .A(Packet_In[13]), .Z(n164) );
  AOI22CDNM1P U77 ( .A(n14), .B(n164), .C(\Queue[4][13] ), .D(n14), .Z(n386)
         );
  N1M1P U78 ( .A(Packet_In[14]), .Z(n166) );
  AOI22CDNM1P U79 ( .A(n14), .B(n166), .C(\Queue[4][14] ), .D(n14), .Z(n387)
         );
  N1M1P U80 ( .A(Packet_In[15]), .Z(n168) );
  AOI22CDNM1P U81 ( .A(n14), .B(n168), .C(\Queue[4][15] ), .D(n14), .Z(n388)
         );
  N1M1P U82 ( .A(Packet_In[16]), .Z(n170) );
  AOI22CDNM1P U83 ( .A(n14), .B(n170), .C(\Queue[4][16] ), .D(n14), .Z(n389)
         );
  N1M1P U84 ( .A(Packet_In[17]), .Z(n172) );
  AOI22CDNM1P U85 ( .A(n14), .B(n172), .C(\Queue[4][17] ), .D(n14), .Z(n390)
         );
  N1M1P U86 ( .A(Packet_In[18]), .Z(n174) );
  AOI22CDNM1P U87 ( .A(n14), .B(n174), .C(\Queue[4][18] ), .D(n14), .Z(n391)
         );
  N1M1P U88 ( .A(Packet_In[19]), .Z(n176) );
  AOI22CDNM1P U89 ( .A(n14), .B(n176), .C(\Queue[4][19] ), .D(n14), .Z(n392)
         );
  N1M1P U90 ( .A(Packet_In[20]), .Z(n178) );
  AOI22CDNM1P U91 ( .A(n14), .B(n178), .C(\Queue[4][20] ), .D(n14), .Z(n393)
         );
  N1M1P U92 ( .A(Packet_In[21]), .Z(n180) );
  AOI22CDNM1P U93 ( .A(n14), .B(n180), .C(\Queue[4][21] ), .D(n14), .Z(n394)
         );
  N1M1P U94 ( .A(Packet_In[22]), .Z(n182) );
  AOI22CDNM1P U95 ( .A(n14), .B(n182), .C(\Queue[4][22] ), .D(n14), .Z(n395)
         );
  N1M1P U96 ( .A(Packet_In[23]), .Z(n184) );
  AOI22CDNM1P U97 ( .A(n14), .B(n184), .C(\Queue[4][23] ), .D(n14), .Z(n396)
         );
  N1M1P U98 ( .A(Packet_In[24]), .Z(n186) );
  AOI22CDNM1P U99 ( .A(n14), .B(n186), .C(\Queue[4][24] ), .D(n14), .Z(n397)
         );
  AOI22CDNM1P U100 ( .A(n14), .B(n188), .C(\Queue[4][25] ), .D(n14), .Z(n398)
         );
  N1M1P U101 ( .A(Packet_In[26]), .Z(n190) );
  AOI22CDNM1P U102 ( .A(n14), .B(n190), .C(\Queue[4][26] ), .D(n14), .Z(n399)
         );
  AOI22CDNM1P U103 ( .A(n14), .B(n192), .C(\Queue[4][27] ), .D(n14), .Z(n400)
         );
  N1M1P U104 ( .A(Packet_In[28]), .Z(n194) );
  AOI22CDNM1P U105 ( .A(n14), .B(n194), .C(\Queue[4][28] ), .D(n14), .Z(n401)
         );
  AOI22CDNM1P U106 ( .A(n14), .B(n196), .C(\Queue[4][29] ), .D(n14), .Z(n402)
         );
  AOI22CDNM1P U107 ( .A(n14), .B(n198), .C(\Queue[4][30] ), .D(n14), .Z(n403)
         );
  OAI22CDNM1P U108 ( .A(n133), .B(n15), .C(n204), .D(Full), .Z(n404) );
  OA21M1P U109 ( .A(n133), .B(n206), .C(Rst_n), .Z(n18) );
  AOI22M1P U110 ( .A(\Queue[2][0] ), .B(n51), .C(\Queue[1][0] ), .D(n4), .Z(
        n19) );
  OAI21M1P U111 ( .A(n138), .B(n53), .C(n19), .Z(n405) );
  AOI22M1P U112 ( .A(n51), .B(\Queue[2][1] ), .C(\Queue[1][1] ), .D(n4), .Z(
        n20) );
  OAI21M1P U113 ( .A(n53), .B(n140), .C(n20), .Z(n406) );
  AOI22M1P U114 ( .A(n51), .B(\Queue[2][2] ), .C(\Queue[1][2] ), .D(n4), .Z(
        n21) );
  OAI21M1P U115 ( .A(n53), .B(n142), .C(n21), .Z(n407) );
  AOI22M1P U116 ( .A(n51), .B(\Queue[2][3] ), .C(\Queue[1][3] ), .D(n4), .Z(
        n22) );
  OAI21M1P U117 ( .A(n53), .B(n144), .C(n22), .Z(n408) );
  AOI22M1P U118 ( .A(n51), .B(\Queue[2][4] ), .C(\Queue[1][4] ), .D(n4), .Z(
        n23) );
  OAI21M1P U119 ( .A(n53), .B(n146), .C(n23), .Z(n409) );
  AOI22M1P U120 ( .A(n51), .B(\Queue[2][5] ), .C(\Queue[1][5] ), .D(n4), .Z(
        n24) );
  OAI21M1P U121 ( .A(n53), .B(n148), .C(n24), .Z(n410) );
  AOI22M1P U122 ( .A(n51), .B(\Queue[2][6] ), .C(\Queue[1][6] ), .D(n4), .Z(
        n25) );
  OAI21M1P U123 ( .A(n53), .B(n150), .C(n25), .Z(n411) );
  AOI22M1P U124 ( .A(n51), .B(\Queue[2][7] ), .C(\Queue[1][7] ), .D(n4), .Z(
        n26) );
  OAI21M1P U125 ( .A(n53), .B(n152), .C(n26), .Z(n412) );
  AOI22M1P U126 ( .A(n51), .B(\Queue[2][8] ), .C(\Queue[1][8] ), .D(n4), .Z(
        n27) );
  OAI21M1P U127 ( .A(n53), .B(n154), .C(n27), .Z(n413) );
  AOI22M1P U128 ( .A(n51), .B(\Queue[2][9] ), .C(\Queue[1][9] ), .D(n5), .Z(
        n28) );
  OAI21M1P U129 ( .A(n53), .B(n156), .C(n28), .Z(n414) );
  AOI22M1P U130 ( .A(n51), .B(\Queue[2][10] ), .C(\Queue[1][10] ), .D(n5), .Z(
        n29) );
  OAI21M1P U131 ( .A(n53), .B(n158), .C(n29), .Z(n415) );
  AOI22M1P U132 ( .A(n51), .B(\Queue[2][11] ), .C(\Queue[1][11] ), .D(n5), .Z(
        n30) );
  OAI21M1P U133 ( .A(n53), .B(n160), .C(n30), .Z(n416) );
  AOI22M1P U134 ( .A(n51), .B(\Queue[2][12] ), .C(\Queue[1][12] ), .D(n5), .Z(
        n31) );
  OAI21M1P U135 ( .A(n53), .B(n162), .C(n31), .Z(n417) );
  AOI22M1P U136 ( .A(n51), .B(\Queue[2][13] ), .C(\Queue[1][13] ), .D(n5), .Z(
        n32) );
  OAI21M1P U137 ( .A(n53), .B(n164), .C(n32), .Z(n418) );
  AOI22M1P U138 ( .A(n51), .B(\Queue[2][14] ), .C(\Queue[1][14] ), .D(n5), .Z(
        n33) );
  OAI21M1P U139 ( .A(n53), .B(n166), .C(n33), .Z(n419) );
  AOI22M1P U140 ( .A(n51), .B(\Queue[2][15] ), .C(\Queue[1][15] ), .D(n5), .Z(
        n34) );
  OAI21M1P U141 ( .A(n53), .B(n168), .C(n34), .Z(n420) );
  AOI22M1P U142 ( .A(n51), .B(\Queue[2][16] ), .C(\Queue[1][16] ), .D(n5), .Z(
        n35) );
  OAI21M1P U143 ( .A(n53), .B(n170), .C(n35), .Z(n421) );
  AOI22M1P U144 ( .A(n51), .B(\Queue[2][17] ), .C(\Queue[1][17] ), .D(n5), .Z(
        n36) );
  OAI21M1P U145 ( .A(n53), .B(n172), .C(n36), .Z(n422) );
  AOI22M1P U146 ( .A(n51), .B(\Queue[2][18] ), .C(\Queue[1][18] ), .D(n50), 
        .Z(n37) );
  OAI21M1P U147 ( .A(n53), .B(n174), .C(n37), .Z(n423) );
  AOI22M1P U148 ( .A(n51), .B(\Queue[2][19] ), .C(\Queue[1][19] ), .D(n50), 
        .Z(n38) );
  OAI21M1P U149 ( .A(n53), .B(n176), .C(n38), .Z(n424) );
  AOI22M1P U150 ( .A(n51), .B(\Queue[2][20] ), .C(\Queue[1][20] ), .D(n50), 
        .Z(n39) );
  OAI21M1P U151 ( .A(n53), .B(n178), .C(n39), .Z(n425) );
  AOI22M1P U152 ( .A(n51), .B(\Queue[2][21] ), .C(\Queue[1][21] ), .D(n50), 
        .Z(n40) );
  OAI21M1P U153 ( .A(n53), .B(n180), .C(n40), .Z(n426) );
  AOI22M1P U154 ( .A(n51), .B(\Queue[2][22] ), .C(\Queue[1][22] ), .D(n50), 
        .Z(n41) );
  OAI21M1P U155 ( .A(n53), .B(n182), .C(n41), .Z(n427) );
  AOI22M1P U156 ( .A(n51), .B(\Queue[2][23] ), .C(\Queue[1][23] ), .D(n50), 
        .Z(n42) );
  OAI21M1P U157 ( .A(n53), .B(n184), .C(n42), .Z(n428) );
  AOI22M1P U158 ( .A(n51), .B(\Queue[2][24] ), .C(\Queue[1][24] ), .D(n50), 
        .Z(n43) );
  OAI21M1P U159 ( .A(n53), .B(n186), .C(n43), .Z(n429) );
  AOI22M1P U160 ( .A(n51), .B(\Queue[2][25] ), .C(\Queue[1][25] ), .D(n50), 
        .Z(n44) );
  OAI21M1P U161 ( .A(n53), .B(n188), .C(n44), .Z(n430) );
  AOI22M1P U162 ( .A(n51), .B(\Queue[2][26] ), .C(\Queue[1][26] ), .D(n5), .Z(
        n45) );
  OAI21M1P U163 ( .A(n53), .B(n190), .C(n45), .Z(n431) );
  AOI22M1P U164 ( .A(n51), .B(\Queue[2][27] ), .C(\Queue[1][27] ), .D(n4), .Z(
        n46) );
  OAI21M1P U165 ( .A(n53), .B(n192), .C(n46), .Z(n432) );
  AOI22M1P U166 ( .A(n51), .B(\Queue[2][28] ), .C(\Queue[1][28] ), .D(n4), .Z(
        n47) );
  OAI21M1P U167 ( .A(n53), .B(n194), .C(n47), .Z(n433) );
  AOI22M1P U168 ( .A(n51), .B(\Queue[2][29] ), .C(\Queue[1][29] ), .D(n4), .Z(
        n48) );
  OAI21M1P U169 ( .A(n53), .B(n196), .C(n48), .Z(n434) );
  AOI22M1P U170 ( .A(n51), .B(\Queue[2][30] ), .C(\Queue[1][30] ), .D(n5), .Z(
        n49) );
  OAI21M1P U171 ( .A(n53), .B(n198), .C(n49), .Z(n435) );
  AOI22M1P U172 ( .A(n51), .B(\Queue[2][31] ), .C(\Queue[1][31] ), .D(n5), .Z(
        n52) );
  OAI21M1P U173 ( .A(n53), .B(n203), .C(n52), .Z(n436) );
  OAI21M1P U174 ( .A(n55), .B(n54), .C(n135), .Z(n56) );
  AOI21M1P U175 ( .A(n3), .B(n206), .C(n135), .Z(n89) );
  AOI22M1P U176 ( .A(\Queue[1][0] ), .B(n6), .C(n88), .D(Packet_Out[0]), .Z(
        n57) );
  OAI21M1P U177 ( .A(n138), .B(n91), .C(n57), .Z(n437) );
  AOI22M1P U178 ( .A(\Queue[1][1] ), .B(n6), .C(n88), .D(Packet_Out[1]), .Z(
        n58) );
  OAI21M1P U179 ( .A(n140), .B(n91), .C(n58), .Z(n438) );
  AOI22M1P U180 ( .A(\Queue[1][2] ), .B(n6), .C(n88), .D(Packet_Out[2]), .Z(
        n59) );
  OAI21M1P U181 ( .A(n142), .B(n91), .C(n59), .Z(n439) );
  AOI22M1P U182 ( .A(\Queue[1][3] ), .B(n6), .C(n88), .D(Packet_Out[3]), .Z(
        n60) );
  OAI21M1P U183 ( .A(n144), .B(n91), .C(n60), .Z(n440) );
  AOI22M1P U184 ( .A(\Queue[1][4] ), .B(n6), .C(n88), .D(Packet_Out[4]), .Z(
        n61) );
  OAI21M1P U185 ( .A(n146), .B(n91), .C(n61), .Z(n441) );
  AOI22M1P U186 ( .A(\Queue[1][5] ), .B(n6), .C(n88), .D(Packet_Out[5]), .Z(
        n62) );
  OAI21M1P U187 ( .A(n148), .B(n91), .C(n62), .Z(n442) );
  AOI22M1P U188 ( .A(\Queue[1][6] ), .B(n6), .C(n88), .D(Packet_Out[6]), .Z(
        n63) );
  OAI21M1P U189 ( .A(n150), .B(n91), .C(n63), .Z(n443) );
  AOI22M1P U190 ( .A(\Queue[1][7] ), .B(n6), .C(n88), .D(Packet_Out[7]), .Z(
        n64) );
  OAI21M1P U191 ( .A(n152), .B(n91), .C(n64), .Z(n444) );
  AOI22M1P U192 ( .A(\Queue[1][8] ), .B(n6), .C(n88), .D(Packet_Out[8]), .Z(
        n65) );
  OAI21M1P U193 ( .A(n154), .B(n91), .C(n65), .Z(n445) );
  AOI22M1P U194 ( .A(\Queue[1][9] ), .B(n6), .C(n88), .D(Packet_Out[9]), .Z(
        n66) );
  OAI21M1P U195 ( .A(n156), .B(n91), .C(n66), .Z(n446) );
  AOI22M1P U196 ( .A(\Queue[1][10] ), .B(n6), .C(n88), .D(Packet_Out[10]), .Z(
        n67) );
  OAI21M1P U197 ( .A(n158), .B(n91), .C(n67), .Z(n447) );
  AOI22M1P U198 ( .A(\Queue[1][11] ), .B(n6), .C(n88), .D(Packet_Out[11]), .Z(
        n68) );
  OAI21M1P U199 ( .A(n160), .B(n91), .C(n68), .Z(n448) );
  AOI22M1P U200 ( .A(\Queue[1][12] ), .B(n6), .C(n88), .D(Packet_Out[12]), .Z(
        n69) );
  OAI21M1P U201 ( .A(n162), .B(n91), .C(n69), .Z(n449) );
  AOI22M1P U202 ( .A(\Queue[1][13] ), .B(n6), .C(n88), .D(Packet_Out[13]), .Z(
        n70) );
  OAI21M1P U203 ( .A(n164), .B(n91), .C(n70), .Z(n450) );
  AOI22M1P U204 ( .A(\Queue[1][14] ), .B(n6), .C(n88), .D(Packet_Out[14]), .Z(
        n71) );
  OAI21M1P U205 ( .A(n166), .B(n91), .C(n71), .Z(n451) );
  AOI22M1P U206 ( .A(\Queue[1][15] ), .B(n6), .C(n88), .D(Packet_Out[15]), .Z(
        n72) );
  OAI21M1P U207 ( .A(n168), .B(n91), .C(n72), .Z(n452) );
  AOI22M1P U208 ( .A(\Queue[1][16] ), .B(n6), .C(n88), .D(Packet_Out[16]), .Z(
        n73) );
  OAI21M1P U209 ( .A(n170), .B(n91), .C(n73), .Z(n453) );
  AOI22M1P U210 ( .A(\Queue[1][17] ), .B(n6), .C(n88), .D(Packet_Out[17]), .Z(
        n74) );
  OAI21M1P U211 ( .A(n172), .B(n91), .C(n74), .Z(n454) );
  AOI22M1P U212 ( .A(\Queue[1][18] ), .B(n6), .C(n88), .D(Packet_Out[18]), .Z(
        n75) );
  OAI21M1P U213 ( .A(n174), .B(n91), .C(n75), .Z(n455) );
  AOI22M1P U214 ( .A(\Queue[1][19] ), .B(n6), .C(n88), .D(Packet_Out[19]), .Z(
        n76) );
  OAI21M1P U215 ( .A(n176), .B(n91), .C(n76), .Z(n456) );
  AOI22M1P U216 ( .A(\Queue[1][20] ), .B(n89), .C(n88), .D(Packet_Out[20]), 
        .Z(n77) );
  OAI21M1P U217 ( .A(n178), .B(n91), .C(n77), .Z(n457) );
  AOI22M1P U218 ( .A(\Queue[1][21] ), .B(n89), .C(n88), .D(Packet_Out[21]), 
        .Z(n78) );
  OAI21M1P U219 ( .A(n180), .B(n91), .C(n78), .Z(n458) );
  AOI22M1P U220 ( .A(\Queue[1][22] ), .B(n89), .C(n88), .D(Packet_Out[22]), 
        .Z(n79) );
  OAI21M1P U221 ( .A(n182), .B(n91), .C(n79), .Z(n459) );
  AOI22M1P U222 ( .A(\Queue[1][23] ), .B(n89), .C(n88), .D(Packet_Out[23]), 
        .Z(n80) );
  OAI21M1P U223 ( .A(n184), .B(n91), .C(n80), .Z(n460) );
  AOI22M1P U224 ( .A(\Queue[1][24] ), .B(n89), .C(n88), .D(Packet_Out[24]), 
        .Z(n81) );
  OAI21M1P U225 ( .A(n186), .B(n91), .C(n81), .Z(n461) );
  AOI22M1P U226 ( .A(\Queue[1][25] ), .B(n89), .C(n88), .D(Packet_Out[25]), 
        .Z(n82) );
  OAI21M1P U227 ( .A(n188), .B(n91), .C(n82), .Z(n462) );
  AOI22M1P U228 ( .A(\Queue[1][26] ), .B(n6), .C(n88), .D(Packet_Out[26]), .Z(
        n83) );
  OAI21M1P U229 ( .A(n190), .B(n91), .C(n83), .Z(n463) );
  AOI22M1P U230 ( .A(\Queue[1][27] ), .B(n6), .C(n88), .D(Packet_Out[27]), .Z(
        n84) );
  OAI21M1P U231 ( .A(n192), .B(n91), .C(n84), .Z(n464) );
  AOI22M1P U232 ( .A(\Queue[1][28] ), .B(n6), .C(n88), .D(Packet_Out[28]), .Z(
        n85) );
  OAI21M1P U233 ( .A(n194), .B(n91), .C(n85), .Z(n465) );
  AOI22M1P U234 ( .A(\Queue[1][29] ), .B(n6), .C(n88), .D(Packet_Out[29]), .Z(
        n86) );
  OAI21M1P U235 ( .A(n196), .B(n91), .C(n86), .Z(n466) );
  AOI22M1P U236 ( .A(\Queue[1][30] ), .B(n6), .C(n88), .D(Packet_Out[30]), .Z(
        n87) );
  OAI21M1P U237 ( .A(n198), .B(n91), .C(n87), .Z(n467) );
  AOI22M1P U238 ( .A(\Queue[1][31] ), .B(n6), .C(n88), .D(Packet_Out[31]), .Z(
        n90) );
  OAI21M1P U239 ( .A(n203), .B(n91), .C(n90), .Z(n468) );
  OA21M1P U240 ( .A(n133), .B(n94), .C(Rst_n), .Z(n92) );
  ND2M1P U241 ( .A(n93), .B(n131), .Z(n132) );
  AOI22M1P U242 ( .A(\Queue[2][0] ), .B(n127), .C(\Queue[3][0] ), .D(n126), 
        .Z(n95) );
  OAI21M1P U243 ( .A(n138), .B(n129), .C(n95), .Z(n469) );
  AOI22M1P U244 ( .A(\Queue[2][1] ), .B(n127), .C(n126), .D(\Queue[3][1] ), 
        .Z(n96) );
  OAI21M1P U245 ( .A(n140), .B(n129), .C(n96), .Z(n470) );
  AOI22M1P U246 ( .A(\Queue[2][2] ), .B(n127), .C(n126), .D(\Queue[3][2] ), 
        .Z(n97) );
  OAI21M1P U247 ( .A(n142), .B(n129), .C(n97), .Z(n471) );
  AOI22M1P U248 ( .A(\Queue[2][3] ), .B(n127), .C(n126), .D(\Queue[3][3] ), 
        .Z(n98) );
  OAI21M1P U249 ( .A(n144), .B(n129), .C(n98), .Z(n472) );
  AOI22M1P U250 ( .A(\Queue[2][4] ), .B(n127), .C(n126), .D(\Queue[3][4] ), 
        .Z(n99) );
  OAI21M1P U251 ( .A(n146), .B(n129), .C(n99), .Z(n473) );
  AOI22M1P U252 ( .A(\Queue[2][5] ), .B(n127), .C(n126), .D(\Queue[3][5] ), 
        .Z(n100) );
  OAI21M1P U253 ( .A(n148), .B(n129), .C(n100), .Z(n474) );
  AOI22M1P U254 ( .A(\Queue[2][6] ), .B(n127), .C(n126), .D(\Queue[3][6] ), 
        .Z(n101) );
  OAI21M1P U255 ( .A(n150), .B(n129), .C(n101), .Z(n475) );
  AOI22M1P U256 ( .A(\Queue[2][7] ), .B(n127), .C(n126), .D(\Queue[3][7] ), 
        .Z(n102) );
  OAI21M1P U257 ( .A(n152), .B(n129), .C(n102), .Z(n476) );
  AOI22M1P U258 ( .A(\Queue[2][8] ), .B(n127), .C(n126), .D(\Queue[3][8] ), 
        .Z(n103) );
  OAI21M1P U259 ( .A(n154), .B(n129), .C(n103), .Z(n477) );
  AOI22M1P U260 ( .A(\Queue[2][9] ), .B(n127), .C(n126), .D(\Queue[3][9] ), 
        .Z(n104) );
  OAI21M1P U261 ( .A(n156), .B(n129), .C(n104), .Z(n478) );
  AOI22M1P U262 ( .A(\Queue[2][10] ), .B(n127), .C(n126), .D(\Queue[3][10] ), 
        .Z(n105) );
  OAI21M1P U263 ( .A(n158), .B(n129), .C(n105), .Z(n479) );
  AOI22M1P U264 ( .A(\Queue[2][11] ), .B(n127), .C(n126), .D(\Queue[3][11] ), 
        .Z(n106) );
  OAI21M1P U265 ( .A(n160), .B(n129), .C(n106), .Z(n480) );
  AOI22M1P U266 ( .A(\Queue[2][12] ), .B(n127), .C(n126), .D(\Queue[3][12] ), 
        .Z(n107) );
  OAI21M1P U267 ( .A(n162), .B(n129), .C(n107), .Z(n481) );
  AOI22M1P U268 ( .A(\Queue[2][13] ), .B(n127), .C(n126), .D(\Queue[3][13] ), 
        .Z(n108) );
  OAI21M1P U269 ( .A(n164), .B(n129), .C(n108), .Z(n482) );
  AOI22M1P U270 ( .A(\Queue[2][14] ), .B(n127), .C(n126), .D(\Queue[3][14] ), 
        .Z(n109) );
  OAI21M1P U271 ( .A(n166), .B(n129), .C(n109), .Z(n483) );
  AOI22M1P U272 ( .A(\Queue[2][15] ), .B(n127), .C(n126), .D(\Queue[3][15] ), 
        .Z(n110) );
  OAI21M1P U273 ( .A(n168), .B(n129), .C(n110), .Z(n484) );
  AOI22M1P U274 ( .A(\Queue[2][16] ), .B(n127), .C(n126), .D(\Queue[3][16] ), 
        .Z(n111) );
  OAI21M1P U275 ( .A(n170), .B(n129), .C(n111), .Z(n485) );
  AOI22M1P U276 ( .A(\Queue[2][17] ), .B(n127), .C(n126), .D(\Queue[3][17] ), 
        .Z(n112) );
  OAI21M1P U277 ( .A(n172), .B(n129), .C(n112), .Z(n486) );
  AOI22M1P U278 ( .A(\Queue[2][18] ), .B(n127), .C(n126), .D(\Queue[3][18] ), 
        .Z(n113) );
  OAI21M1P U279 ( .A(n174), .B(n129), .C(n113), .Z(n487) );
  AOI22M1P U280 ( .A(\Queue[2][19] ), .B(n127), .C(n126), .D(\Queue[3][19] ), 
        .Z(n114) );
  OAI21M1P U281 ( .A(n176), .B(n129), .C(n114), .Z(n488) );
  AOI22M1P U282 ( .A(\Queue[2][20] ), .B(n127), .C(n126), .D(\Queue[3][20] ), 
        .Z(n115) );
  OAI21M1P U283 ( .A(n178), .B(n129), .C(n115), .Z(n489) );
  AOI22M1P U284 ( .A(\Queue[2][21] ), .B(n127), .C(n126), .D(\Queue[3][21] ), 
        .Z(n116) );
  OAI21M1P U285 ( .A(n180), .B(n129), .C(n116), .Z(n490) );
  AOI22M1P U286 ( .A(\Queue[2][22] ), .B(n127), .C(n126), .D(\Queue[3][22] ), 
        .Z(n117) );
  OAI21M1P U287 ( .A(n182), .B(n129), .C(n117), .Z(n491) );
  AOI22M1P U288 ( .A(\Queue[2][23] ), .B(n127), .C(n126), .D(\Queue[3][23] ), 
        .Z(n118) );
  OAI21M1P U289 ( .A(n184), .B(n129), .C(n118), .Z(n492) );
  AOI22M1P U290 ( .A(\Queue[2][24] ), .B(n127), .C(n126), .D(\Queue[3][24] ), 
        .Z(n119) );
  OAI21M1P U291 ( .A(n186), .B(n129), .C(n119), .Z(n493) );
  AOI22M1P U292 ( .A(\Queue[2][25] ), .B(n127), .C(n126), .D(\Queue[3][25] ), 
        .Z(n120) );
  OAI21M1P U293 ( .A(n188), .B(n129), .C(n120), .Z(n494) );
  AOI22M1P U294 ( .A(\Queue[2][26] ), .B(n127), .C(n126), .D(\Queue[3][26] ), 
        .Z(n121) );
  OAI21M1P U295 ( .A(n190), .B(n129), .C(n121), .Z(n495) );
  AOI22M1P U296 ( .A(\Queue[2][27] ), .B(n127), .C(n126), .D(\Queue[3][27] ), 
        .Z(n122) );
  OAI21M1P U297 ( .A(n192), .B(n129), .C(n122), .Z(n496) );
  AOI22M1P U298 ( .A(\Queue[2][28] ), .B(n127), .C(n126), .D(\Queue[3][28] ), 
        .Z(n123) );
  OAI21M1P U299 ( .A(n194), .B(n129), .C(n123), .Z(n497) );
  AOI22M1P U300 ( .A(\Queue[2][29] ), .B(n127), .C(n126), .D(\Queue[3][29] ), 
        .Z(n124) );
  OAI21M1P U301 ( .A(n196), .B(n129), .C(n124), .Z(n498) );
  AOI22M1P U302 ( .A(\Queue[2][30] ), .B(n127), .C(n126), .D(\Queue[3][30] ), 
        .Z(n125) );
  OAI21M1P U303 ( .A(n198), .B(n129), .C(n125), .Z(n499) );
  AOI22M1P U304 ( .A(\Queue[2][31] ), .B(n127), .C(n126), .D(\Queue[3][31] ), 
        .Z(n128) );
  OAI21M1P U305 ( .A(n203), .B(n129), .C(n128), .Z(n500) );
  OA21M1P U306 ( .A(n133), .B(n134), .C(Rst_n), .Z(n130) );
  AOI22M1P U307 ( .A(\Queue[3][0] ), .B(n200), .C(n199), .D(\Queue[4][0] ), 
        .Z(n137) );
  OAI21M1P U308 ( .A(n138), .B(n202), .C(n137), .Z(n501) );
  AOI22M1P U309 ( .A(\Queue[3][1] ), .B(n200), .C(n199), .D(\Queue[4][1] ), 
        .Z(n139) );
  OAI21M1P U310 ( .A(n140), .B(n202), .C(n139), .Z(n502) );
  AOI22M1P U311 ( .A(\Queue[3][2] ), .B(n200), .C(n199), .D(\Queue[4][2] ), 
        .Z(n141) );
  OAI21M1P U312 ( .A(n142), .B(n202), .C(n141), .Z(n503) );
  AOI22M1P U313 ( .A(\Queue[3][3] ), .B(n200), .C(n199), .D(\Queue[4][3] ), 
        .Z(n143) );
  OAI21M1P U314 ( .A(n144), .B(n202), .C(n143), .Z(n504) );
  AOI22M1P U315 ( .A(\Queue[3][4] ), .B(n200), .C(n199), .D(\Queue[4][4] ), 
        .Z(n145) );
  OAI21M1P U316 ( .A(n146), .B(n202), .C(n145), .Z(n505) );
  AOI22M1P U317 ( .A(\Queue[3][5] ), .B(n200), .C(n199), .D(\Queue[4][5] ), 
        .Z(n147) );
  OAI21M1P U318 ( .A(n148), .B(n202), .C(n147), .Z(n506) );
  AOI22M1P U319 ( .A(\Queue[3][6] ), .B(n200), .C(n199), .D(\Queue[4][6] ), 
        .Z(n149) );
  OAI21M1P U320 ( .A(n150), .B(n202), .C(n149), .Z(n507) );
  AOI22M1P U321 ( .A(\Queue[3][7] ), .B(n200), .C(n199), .D(\Queue[4][7] ), 
        .Z(n151) );
  OAI21M1P U322 ( .A(n152), .B(n202), .C(n151), .Z(n508) );
  AOI22M1P U323 ( .A(\Queue[3][8] ), .B(n200), .C(n199), .D(\Queue[4][8] ), 
        .Z(n153) );
  OAI21M1P U324 ( .A(n154), .B(n202), .C(n153), .Z(n509) );
  AOI22M1P U325 ( .A(\Queue[3][9] ), .B(n200), .C(n199), .D(\Queue[4][9] ), 
        .Z(n155) );
  OAI21M1P U326 ( .A(n156), .B(n202), .C(n155), .Z(n510) );
  AOI22M1P U327 ( .A(\Queue[3][10] ), .B(n200), .C(n199), .D(\Queue[4][10] ), 
        .Z(n157) );
  OAI21M1P U328 ( .A(n158), .B(n202), .C(n157), .Z(n511) );
  AOI22M1P U329 ( .A(\Queue[3][11] ), .B(n200), .C(n199), .D(\Queue[4][11] ), 
        .Z(n159) );
  OAI21M1P U330 ( .A(n160), .B(n202), .C(n159), .Z(n512) );
  AOI22M1P U331 ( .A(\Queue[3][12] ), .B(n200), .C(n199), .D(\Queue[4][12] ), 
        .Z(n161) );
  OAI21M1P U332 ( .A(n162), .B(n202), .C(n161), .Z(n513) );
  AOI22M1P U333 ( .A(\Queue[3][13] ), .B(n200), .C(n199), .D(\Queue[4][13] ), 
        .Z(n163) );
  OAI21M1P U334 ( .A(n164), .B(n202), .C(n163), .Z(n514) );
  AOI22M1P U335 ( .A(\Queue[3][14] ), .B(n200), .C(n199), .D(\Queue[4][14] ), 
        .Z(n165) );
  OAI21M1P U336 ( .A(n166), .B(n202), .C(n165), .Z(n515) );
  AOI22M1P U337 ( .A(\Queue[3][15] ), .B(n200), .C(n199), .D(\Queue[4][15] ), 
        .Z(n167) );
  OAI21M1P U338 ( .A(n168), .B(n202), .C(n167), .Z(n516) );
  AOI22M1P U339 ( .A(\Queue[3][16] ), .B(n200), .C(n199), .D(\Queue[4][16] ), 
        .Z(n169) );
  OAI21M1P U340 ( .A(n170), .B(n202), .C(n169), .Z(n517) );
  AOI22M1P U341 ( .A(\Queue[3][17] ), .B(n200), .C(n199), .D(\Queue[4][17] ), 
        .Z(n171) );
  OAI21M1P U342 ( .A(n172), .B(n202), .C(n171), .Z(n518) );
  AOI22M1P U343 ( .A(\Queue[3][18] ), .B(n200), .C(n199), .D(\Queue[4][18] ), 
        .Z(n173) );
  OAI21M1P U344 ( .A(n174), .B(n202), .C(n173), .Z(n519) );
  AOI22M1P U345 ( .A(\Queue[3][19] ), .B(n200), .C(n199), .D(\Queue[4][19] ), 
        .Z(n175) );
  OAI21M1P U346 ( .A(n176), .B(n202), .C(n175), .Z(n520) );
  AOI22M1P U347 ( .A(\Queue[3][20] ), .B(n200), .C(n199), .D(\Queue[4][20] ), 
        .Z(n177) );
  OAI21M1P U348 ( .A(n178), .B(n202), .C(n177), .Z(n521) );
  AOI22M1P U349 ( .A(\Queue[3][21] ), .B(n200), .C(n199), .D(\Queue[4][21] ), 
        .Z(n179) );
  OAI21M1P U350 ( .A(n180), .B(n202), .C(n179), .Z(n522) );
  AOI22M1P U351 ( .A(\Queue[3][22] ), .B(n200), .C(n199), .D(\Queue[4][22] ), 
        .Z(n181) );
  OAI21M1P U352 ( .A(n182), .B(n202), .C(n181), .Z(n523) );
  AOI22M1P U353 ( .A(\Queue[3][23] ), .B(n200), .C(n199), .D(\Queue[4][23] ), 
        .Z(n183) );
  OAI21M1P U354 ( .A(n184), .B(n202), .C(n183), .Z(n524) );
  AOI22M1P U355 ( .A(\Queue[3][24] ), .B(n200), .C(n199), .D(\Queue[4][24] ), 
        .Z(n185) );
  OAI21M1P U356 ( .A(n186), .B(n202), .C(n185), .Z(n525) );
  AOI22M1P U357 ( .A(\Queue[3][25] ), .B(n200), .C(n199), .D(\Queue[4][25] ), 
        .Z(n187) );
  OAI21M1P U358 ( .A(n188), .B(n202), .C(n187), .Z(n526) );
  AOI22M1P U359 ( .A(\Queue[3][26] ), .B(n200), .C(n199), .D(\Queue[4][26] ), 
        .Z(n189) );
  OAI21M1P U360 ( .A(n190), .B(n202), .C(n189), .Z(n527) );
  AOI22M1P U361 ( .A(\Queue[3][27] ), .B(n200), .C(n199), .D(\Queue[4][27] ), 
        .Z(n191) );
  OAI21M1P U362 ( .A(n192), .B(n202), .C(n191), .Z(n528) );
  AOI22M1P U363 ( .A(\Queue[3][28] ), .B(n200), .C(n199), .D(\Queue[4][28] ), 
        .Z(n193) );
  OAI21M1P U364 ( .A(n194), .B(n202), .C(n193), .Z(n529) );
  AOI22M1P U365 ( .A(\Queue[3][29] ), .B(n200), .C(n199), .D(\Queue[4][29] ), 
        .Z(n195) );
  OAI21M1P U366 ( .A(n196), .B(n202), .C(n195), .Z(n530) );
  AOI22M1P U367 ( .A(\Queue[3][30] ), .B(n200), .C(n199), .D(\Queue[4][30] ), 
        .Z(n197) );
  OAI21M1P U368 ( .A(n198), .B(n202), .C(n197), .Z(n531) );
  AOI22M1P U369 ( .A(\Queue[3][31] ), .B(n200), .C(n199), .D(\Queue[4][31] ), 
        .Z(n201) );
  OAI21M1P U370 ( .A(n203), .B(n202), .C(n201), .Z(n532) );
  N1M1P U371 ( .A(n533), .Z(Empty) );
  AOI22M1P U372 ( .A(n206), .B(n205), .C(n204), .D(Empty), .Z(n534) );
endmodule


module Packet_Queue_2 ( Clk_r, Rst_n, Packet_In, Read_Ack, Write_Ack, 
        Packet_Out, Empty, Full );
  input [31:0] Packet_In;
  output [31:0] Packet_Out;
  input Clk_r, Rst_n, Read_Ack, Write_Ack;
  output Empty, Full;
  wire   \Queue[4][31] , \Queue[4][30] , \Queue[4][29] , \Queue[4][28] ,
         \Queue[4][27] , \Queue[4][26] , \Queue[4][25] , \Queue[4][24] ,
         \Queue[4][15] , \Queue[4][14] , \Queue[4][13] , \Queue[4][12] ,
         \Queue[4][11] , \Queue[4][10] , \Queue[4][9] , \Queue[4][8] ,
         \Queue[4][7] , \Queue[4][6] , \Queue[4][5] , \Queue[4][4] ,
         \Queue[4][3] , \Queue[4][2] , \Queue[4][1] , \Queue[4][0] ,
         \Queue[3][31] , \Queue[3][30] , \Queue[3][29] , \Queue[3][28] ,
         \Queue[3][27] , \Queue[3][26] , \Queue[3][25] , \Queue[3][24] ,
         \Queue[3][15] , \Queue[3][14] , \Queue[3][13] , \Queue[3][12] ,
         \Queue[3][11] , \Queue[3][10] , \Queue[3][9] , \Queue[3][8] ,
         \Queue[3][7] , \Queue[3][6] , \Queue[3][5] , \Queue[3][4] ,
         \Queue[3][3] , \Queue[3][2] , \Queue[3][1] , \Queue[3][0] ,
         \Queue[2][31] , \Queue[2][30] , \Queue[2][29] , \Queue[2][28] ,
         \Queue[2][27] , \Queue[2][26] , \Queue[2][25] , \Queue[2][24] ,
         \Queue[2][15] , \Queue[2][14] , \Queue[2][13] , \Queue[2][12] ,
         \Queue[2][11] , \Queue[2][10] , \Queue[2][9] , \Queue[2][8] ,
         \Queue[2][7] , \Queue[2][6] , \Queue[2][5] , \Queue[2][4] ,
         \Queue[2][3] , \Queue[2][2] , \Queue[2][1] , \Queue[2][0] ,
         \Queue[1][31] , \Queue[1][30] , \Queue[1][29] , \Queue[1][28] ,
         \Queue[1][27] , \Queue[1][26] , \Queue[1][25] , \Queue[1][24] ,
         \Queue[1][15] , \Queue[1][14] , \Queue[1][13] , \Queue[1][12] ,
         \Queue[1][11] , \Queue[1][10] , \Queue[1][9] , \Queue[1][8] ,
         \Queue[1][7] , \Queue[1][6] , \Queue[1][5] , \Queue[1][4] ,
         \Queue[1][3] , \Queue[1][2] , \Queue[1][1] , \Queue[1][0] , n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n217, n218, n219, n220,
         n221, n222, n223, n224, n249, n250, n251, n252, n253, n254, n255,
         n256, n281, n282, n283, n284, n285, n286, n287, n288, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356;
  wire   [2:0] Count;

  FDN2QM1P \Count_reg[0]  ( .D(n170), .CPN(Clk_r), .CD(Rst_n), .Q(Count[0]) );
  FDN2QM1P \Count_reg[1]  ( .D(n171), .CPN(Clk_r), .CD(Rst_n), .Q(Count[1]) );
  FDN2QM1P \Count_reg[2]  ( .D(n172), .CPN(Clk_r), .CD(Rst_n), .Q(Count[2]) );
  FDN1QM1P \Queue_reg[4][30]  ( .D(n196), .CPN(Clk_r), .Q(\Queue[4][30] ) );
  FDN1QM1P \Queue_reg[3][30]  ( .D(n353), .CPN(Clk_r), .Q(\Queue[3][30] ) );
  FDN1QM1P \Queue_reg[2][30]  ( .D(n329), .CPN(Clk_r), .Q(\Queue[2][30] ) );
  FDN1QM1P \Queue_reg[4][29]  ( .D(n195), .CPN(Clk_r), .Q(\Queue[4][29] ) );
  FDN1QM1P \Queue_reg[3][29]  ( .D(n352), .CPN(Clk_r), .Q(\Queue[3][29] ) );
  FDN1QM1P \Queue_reg[2][29]  ( .D(n328), .CPN(Clk_r), .Q(\Queue[2][29] ) );
  FDN1QM1P \Queue_reg[4][28]  ( .D(n194), .CPN(Clk_r), .Q(\Queue[4][28] ) );
  FDN1QM1P \Queue_reg[3][28]  ( .D(n351), .CPN(Clk_r), .Q(\Queue[3][28] ) );
  FDN1QM1P \Queue_reg[2][28]  ( .D(n327), .CPN(Clk_r), .Q(\Queue[2][28] ) );
  FDN1QM1P \Queue_reg[4][27]  ( .D(n193), .CPN(Clk_r), .Q(\Queue[4][27] ) );
  FDN1QM1P \Queue_reg[3][27]  ( .D(n350), .CPN(Clk_r), .Q(\Queue[3][27] ) );
  FDN1QM1P \Queue_reg[2][27]  ( .D(n326), .CPN(Clk_r), .Q(\Queue[2][27] ) );
  FDN1QM1P \Queue_reg[4][26]  ( .D(n192), .CPN(Clk_r), .Q(\Queue[4][26] ) );
  FDN1QM1P \Queue_reg[3][26]  ( .D(n349), .CPN(Clk_r), .Q(\Queue[3][26] ) );
  FDN1QM1P \Queue_reg[2][26]  ( .D(n325), .CPN(Clk_r), .Q(\Queue[2][26] ) );
  FDN1QM1P \Queue_reg[4][25]  ( .D(n191), .CPN(Clk_r), .Q(\Queue[4][25] ) );
  FDN1QM1P \Queue_reg[3][25]  ( .D(n348), .CPN(Clk_r), .Q(\Queue[3][25] ) );
  FDN1QM1P \Queue_reg[2][25]  ( .D(n324), .CPN(Clk_r), .Q(\Queue[2][25] ) );
  FDN1QM1P \Queue_reg[4][24]  ( .D(n190), .CPN(Clk_r), .Q(\Queue[4][24] ) );
  FDN1QM1P \Queue_reg[3][24]  ( .D(n347), .CPN(Clk_r), .Q(\Queue[3][24] ) );
  FDN1QM1P \Queue_reg[2][24]  ( .D(n323), .CPN(Clk_r), .Q(\Queue[2][24] ) );
  FDN1QM1P \Queue_reg[4][15]  ( .D(n189), .CPN(Clk_r), .Q(\Queue[4][15] ) );
  FDN1QM1P \Queue_reg[3][15]  ( .D(n346), .CPN(Clk_r), .Q(\Queue[3][15] ) );
  FDN1QM1P \Queue_reg[2][15]  ( .D(n322), .CPN(Clk_r), .Q(\Queue[2][15] ) );
  FDN1QM1P \Queue_reg[4][14]  ( .D(n188), .CPN(Clk_r), .Q(\Queue[4][14] ) );
  FDN1QM1P \Queue_reg[3][14]  ( .D(n345), .CPN(Clk_r), .Q(\Queue[3][14] ) );
  FDN1QM1P \Queue_reg[2][14]  ( .D(n321), .CPN(Clk_r), .Q(\Queue[2][14] ) );
  FDN1QM1P \Queue_reg[4][13]  ( .D(n187), .CPN(Clk_r), .Q(\Queue[4][13] ) );
  FDN1QM1P \Queue_reg[3][13]  ( .D(n344), .CPN(Clk_r), .Q(\Queue[3][13] ) );
  FDN1QM1P \Queue_reg[2][13]  ( .D(n320), .CPN(Clk_r), .Q(\Queue[2][13] ) );
  FDN1QM1P \Queue_reg[4][12]  ( .D(n186), .CPN(Clk_r), .Q(\Queue[4][12] ) );
  FDN1QM1P \Queue_reg[3][12]  ( .D(n343), .CPN(Clk_r), .Q(\Queue[3][12] ) );
  FDN1QM1P \Queue_reg[2][12]  ( .D(n319), .CPN(Clk_r), .Q(\Queue[2][12] ) );
  FDN1QM1P \Queue_reg[4][11]  ( .D(n185), .CPN(Clk_r), .Q(\Queue[4][11] ) );
  FDN1QM1P \Queue_reg[3][11]  ( .D(n342), .CPN(Clk_r), .Q(\Queue[3][11] ) );
  FDN1QM1P \Queue_reg[2][11]  ( .D(n318), .CPN(Clk_r), .Q(\Queue[2][11] ) );
  FDN1QM1P \Queue_reg[4][10]  ( .D(n184), .CPN(Clk_r), .Q(\Queue[4][10] ) );
  FDN1QM1P \Queue_reg[3][10]  ( .D(n341), .CPN(Clk_r), .Q(\Queue[3][10] ) );
  FDN1QM1P \Queue_reg[2][10]  ( .D(n317), .CPN(Clk_r), .Q(\Queue[2][10] ) );
  FDN1QM1P \Queue_reg[4][9]  ( .D(n183), .CPN(Clk_r), .Q(\Queue[4][9] ) );
  FDN1QM1P \Queue_reg[3][9]  ( .D(n340), .CPN(Clk_r), .Q(\Queue[3][9] ) );
  FDN1QM1P \Queue_reg[2][9]  ( .D(n316), .CPN(Clk_r), .Q(\Queue[2][9] ) );
  FDN1QM1P \Queue_reg[4][8]  ( .D(n182), .CPN(Clk_r), .Q(\Queue[4][8] ) );
  FDN1QM1P \Queue_reg[3][8]  ( .D(n339), .CPN(Clk_r), .Q(\Queue[3][8] ) );
  FDN1QM1P \Queue_reg[2][8]  ( .D(n315), .CPN(Clk_r), .Q(\Queue[2][8] ) );
  FDN1QM1P \Queue_reg[4][7]  ( .D(n181), .CPN(Clk_r), .Q(\Queue[4][7] ) );
  FDN1QM1P \Queue_reg[3][7]  ( .D(n338), .CPN(Clk_r), .Q(\Queue[3][7] ) );
  FDN1QM1P \Queue_reg[2][7]  ( .D(n314), .CPN(Clk_r), .Q(\Queue[2][7] ) );
  FDN1QM1P \Queue_reg[4][6]  ( .D(n180), .CPN(Clk_r), .Q(\Queue[4][6] ) );
  FDN1QM1P \Queue_reg[3][6]  ( .D(n337), .CPN(Clk_r), .Q(\Queue[3][6] ) );
  FDN1QM1P \Queue_reg[2][6]  ( .D(n313), .CPN(Clk_r), .Q(\Queue[2][6] ) );
  FDN1QM1P \Queue_reg[4][5]  ( .D(n179), .CPN(Clk_r), .Q(\Queue[4][5] ) );
  FDN1QM1P \Queue_reg[3][5]  ( .D(n336), .CPN(Clk_r), .Q(\Queue[3][5] ) );
  FDN1QM1P \Queue_reg[2][5]  ( .D(n312), .CPN(Clk_r), .Q(\Queue[2][5] ) );
  FDN1QM1P \Queue_reg[4][4]  ( .D(n178), .CPN(Clk_r), .Q(\Queue[4][4] ) );
  FDN1QM1P \Queue_reg[3][4]  ( .D(n335), .CPN(Clk_r), .Q(\Queue[3][4] ) );
  FDN1QM1P \Queue_reg[2][4]  ( .D(n311), .CPN(Clk_r), .Q(\Queue[2][4] ) );
  FDN1QM1P \Queue_reg[4][3]  ( .D(n177), .CPN(Clk_r), .Q(\Queue[4][3] ) );
  FDN1QM1P \Queue_reg[3][3]  ( .D(n334), .CPN(Clk_r), .Q(\Queue[3][3] ) );
  FDN1QM1P \Queue_reg[2][3]  ( .D(n310), .CPN(Clk_r), .Q(\Queue[2][3] ) );
  FDN1QM1P \Queue_reg[4][2]  ( .D(n176), .CPN(Clk_r), .Q(\Queue[4][2] ) );
  FDN1QM1P \Queue_reg[3][2]  ( .D(n333), .CPN(Clk_r), .Q(\Queue[3][2] ) );
  FDN1QM1P \Queue_reg[2][2]  ( .D(n309), .CPN(Clk_r), .Q(\Queue[2][2] ) );
  FDN1QM1P \Queue_reg[4][1]  ( .D(n175), .CPN(Clk_r), .Q(\Queue[4][1] ) );
  FDN1QM1P \Queue_reg[3][1]  ( .D(n332), .CPN(Clk_r), .Q(\Queue[3][1] ) );
  FDN1QM1P \Queue_reg[2][1]  ( .D(n308), .CPN(Clk_r), .Q(\Queue[2][1] ) );
  FDN1QM1P \Queue_reg[4][0]  ( .D(n174), .CPN(Clk_r), .Q(\Queue[4][0] ) );
  FDN1QM1P \Queue_reg[3][0]  ( .D(n331), .CPN(Clk_r), .Q(\Queue[3][0] ) );
  FDN1QM1P \Queue_reg[2][0]  ( .D(n307), .CPN(Clk_r), .Q(\Queue[2][0] ) );
  FDN1QM1P \Queue_reg[4][31]  ( .D(n173), .CPN(Clk_r), .Q(\Queue[4][31] ) );
  FDN1QM1P \Queue_reg[3][31]  ( .D(n354), .CPN(Clk_r), .Q(\Queue[3][31] ) );
  FDN1QM1P \Queue_reg[2][31]  ( .D(n330), .CPN(Clk_r), .Q(\Queue[2][31] ) );
  FDN2QM1P Full_reg ( .D(n197), .CPN(Clk_r), .CD(Rst_n), .Q(Full) );
  FDN1QM1P \Queue_reg[1][31]  ( .D(n253), .CPN(Clk_r), .Q(\Queue[1][31] ) );
  FDN1QM1P \Queue_reg[0][31]  ( .D(n306), .CPN(Clk_r), .Q(Packet_Out[31]) );
  FDN1QM1P \Queue_reg[1][30]  ( .D(n252), .CPN(Clk_r), .Q(\Queue[1][30] ) );
  FDN1QM1P \Queue_reg[0][30]  ( .D(n305), .CPN(Clk_r), .Q(Packet_Out[30]) );
  FDN1QM1P \Queue_reg[1][29]  ( .D(n251), .CPN(Clk_r), .Q(\Queue[1][29] ) );
  FDN1QM1P \Queue_reg[0][29]  ( .D(n304), .CPN(Clk_r), .Q(Packet_Out[29]) );
  FDN1QM1P \Queue_reg[1][28]  ( .D(n250), .CPN(Clk_r), .Q(\Queue[1][28] ) );
  FDN1QM1P \Queue_reg[0][28]  ( .D(n303), .CPN(Clk_r), .Q(Packet_Out[28]) );
  FDN1QM1P \Queue_reg[1][27]  ( .D(n249), .CPN(Clk_r), .Q(\Queue[1][27] ) );
  FDN1QM1P \Queue_reg[0][27]  ( .D(n302), .CPN(Clk_r), .Q(Packet_Out[27]) );
  FDN1QM1P \Queue_reg[1][26]  ( .D(n224), .CPN(Clk_r), .Q(\Queue[1][26] ) );
  FDN1QM1P \Queue_reg[0][26]  ( .D(n301), .CPN(Clk_r), .Q(Packet_Out[26]) );
  FDN1QM1P \Queue_reg[1][25]  ( .D(n223), .CPN(Clk_r), .Q(\Queue[1][25] ) );
  FDN1QM1P \Queue_reg[0][25]  ( .D(n300), .CPN(Clk_r), .Q(Packet_Out[25]) );
  FDN1QM1P \Queue_reg[1][24]  ( .D(n222), .CPN(Clk_r), .Q(\Queue[1][24] ) );
  FDN1QM1P \Queue_reg[0][24]  ( .D(n299), .CPN(Clk_r), .Q(Packet_Out[24]) );
  FDN1QM1P \Queue_reg[1][15]  ( .D(n221), .CPN(Clk_r), .Q(\Queue[1][15] ) );
  FDN1QM1P \Queue_reg[0][15]  ( .D(n298), .CPN(Clk_r), .Q(Packet_Out[15]) );
  FDN1QM1P \Queue_reg[1][14]  ( .D(n220), .CPN(Clk_r), .Q(\Queue[1][14] ) );
  FDN1QM1P \Queue_reg[0][14]  ( .D(n297), .CPN(Clk_r), .Q(Packet_Out[14]) );
  FDN1QM1P \Queue_reg[1][13]  ( .D(n219), .CPN(Clk_r), .Q(\Queue[1][13] ) );
  FDN1QM1P \Queue_reg[0][13]  ( .D(n296), .CPN(Clk_r), .Q(Packet_Out[13]) );
  FDN1QM1P \Queue_reg[1][12]  ( .D(n218), .CPN(Clk_r), .Q(\Queue[1][12] ) );
  FDN1QM1P \Queue_reg[0][12]  ( .D(n295), .CPN(Clk_r), .Q(Packet_Out[12]) );
  FDN1QM1P \Queue_reg[1][11]  ( .D(n217), .CPN(Clk_r), .Q(\Queue[1][11] ) );
  FDN1QM1P \Queue_reg[0][11]  ( .D(n294), .CPN(Clk_r), .Q(Packet_Out[11]) );
  FDN1QM1P \Queue_reg[1][10]  ( .D(n208), .CPN(Clk_r), .Q(\Queue[1][10] ) );
  FDN1QM1P \Queue_reg[0][10]  ( .D(n288), .CPN(Clk_r), .Q(Packet_Out[10]) );
  FDN1QM1P \Queue_reg[1][9]  ( .D(n207), .CPN(Clk_r), .Q(\Queue[1][9] ) );
  FDN1QM1P \Queue_reg[0][9]  ( .D(n287), .CPN(Clk_r), .Q(Packet_Out[9]) );
  FDN1QM1P \Queue_reg[1][8]  ( .D(n206), .CPN(Clk_r), .Q(\Queue[1][8] ) );
  FDN1QM1P \Queue_reg[0][8]  ( .D(n286), .CPN(Clk_r), .Q(Packet_Out[8]) );
  FDN1QM1P \Queue_reg[1][7]  ( .D(n205), .CPN(Clk_r), .Q(\Queue[1][7] ) );
  FDN1QM1P \Queue_reg[0][7]  ( .D(n285), .CPN(Clk_r), .Q(Packet_Out[7]) );
  FDN1QM1P \Queue_reg[1][6]  ( .D(n204), .CPN(Clk_r), .Q(\Queue[1][6] ) );
  FDN1QM1P \Queue_reg[0][6]  ( .D(n284), .CPN(Clk_r), .Q(Packet_Out[6]) );
  FDN1QM1P \Queue_reg[1][5]  ( .D(n203), .CPN(Clk_r), .Q(\Queue[1][5] ) );
  FDN1QM1P \Queue_reg[0][5]  ( .D(n283), .CPN(Clk_r), .Q(Packet_Out[5]) );
  FDN1QM1P \Queue_reg[1][4]  ( .D(n202), .CPN(Clk_r), .Q(\Queue[1][4] ) );
  FDN1QM1P \Queue_reg[0][4]  ( .D(n282), .CPN(Clk_r), .Q(Packet_Out[4]) );
  FDN1QM1P \Queue_reg[1][3]  ( .D(n201), .CPN(Clk_r), .Q(\Queue[1][3] ) );
  FDN1QM1P \Queue_reg[0][3]  ( .D(n281), .CPN(Clk_r), .Q(Packet_Out[3]) );
  FDN1QM1P \Queue_reg[1][2]  ( .D(n200), .CPN(Clk_r), .Q(\Queue[1][2] ) );
  FDN1QM1P \Queue_reg[0][2]  ( .D(n256), .CPN(Clk_r), .Q(Packet_Out[2]) );
  FDN1QM1P \Queue_reg[1][1]  ( .D(n199), .CPN(Clk_r), .Q(\Queue[1][1] ) );
  FDN1QM1P \Queue_reg[0][1]  ( .D(n255), .CPN(Clk_r), .Q(Packet_Out[1]) );
  FDN1QM1P \Queue_reg[1][0]  ( .D(n198), .CPN(Clk_r), .Q(\Queue[1][0] ) );
  FDN1QM1P \Queue_reg[0][0]  ( .D(n254), .CPN(Clk_r), .Q(Packet_Out[0]) );
  FDN2QM1P Empty_reg ( .D(n356), .CPN(Clk_r), .CD(Rst_n), .Q(n355) );
  ND2M1P U3 ( .A(n15), .B(Rst_n), .Z(n50) );
  BUFM2P U4 ( .A(n76), .Z(n4) );
  BUFM2P U5 ( .A(n46), .Z(n6) );
  BUFM2P U6 ( .A(n163), .Z(n9) );
  BUFM2P U7 ( .A(n105), .Z(n5) );
  OAI211M4P U8 ( .A(n115), .B(n110), .C(n7), .D(n109), .Z(n165) );
  NR2FM2P U9 ( .A(n50), .B(n18), .Z(n17) );
  NR3M1P U10 ( .A(Count[0]), .B(Count[2]), .C(n19), .Z(n81) );
  NR3M1P U11 ( .A(n20), .B(Count[2]), .C(Count[1]), .Z(n169) );
  N1M1P U12 ( .A(Read_Ack), .Z(n110) );
  NR3M1P U13 ( .A(Count[2]), .B(n20), .C(n19), .Z(n113) );
  OAI211M4P U14 ( .A(n81), .B(n110), .C(n7), .D(n21), .Z(n48) );
  OAI211M4P U15 ( .A(n113), .B(n110), .C(n7), .D(n79), .Z(n108) );
  OAI211M4P U16 ( .A(n169), .B(n110), .C(n7), .D(n51), .Z(n78) );
  OAI211M4P U17 ( .A(n81), .B(n112), .C(Rst_n), .D(n111), .Z(n106) );
  N1M2P U18 ( .A(n51), .Z(n75) );
  AOI21M2P U19 ( .A(n7), .B(n115), .C(n114), .Z(n162) );
  OAI21M2P U20 ( .A(n7), .B(Read_Ack), .C(n21), .Z(n45) );
  BUFM2P U21 ( .A(n45), .Z(n3) );
  NR3M1P U22 ( .A(Count[0]), .B(Count[1]), .C(n16), .Z(n115) );
  N1M1P U23 ( .A(n115), .Z(n18) );
  N1M1P U24 ( .A(Count[1]), .Z(n19) );
  N1M1P U25 ( .A(Count[0]), .Z(n20) );
  N1M1P U26 ( .A(Count[2]), .Z(n16) );
  ND2M2P U27 ( .A(Read_Ack), .B(Rst_n), .Z(n114) );
  NR2M3P U28 ( .A(Read_Ack), .B(n80), .Z(n15) );
  BUFM3P U29 ( .A(Write_Ack), .Z(n7) );
  N1M1P U30 ( .A(Packet_In[2]), .Z(n121) );
  N1M1P U31 ( .A(Packet_In[0]), .Z(n117) );
  N1M1P U32 ( .A(Packet_In[28]), .Z(n157) );
  N1M1P U33 ( .A(Packet_In[30]), .Z(n161) );
  N1M1P U34 ( .A(Packet_In[31]), .Z(n166) );
  N1M1P U35 ( .A(Packet_In[29]), .Z(n159) );
  N1M1P U36 ( .A(Packet_In[3]), .Z(n123) );
  N1M1P U37 ( .A(Packet_In[13]), .Z(n143) );
  N1M1P U38 ( .A(Packet_In[27]), .Z(n155) );
  N1M1P U39 ( .A(Packet_In[8]), .Z(n133) );
  N1M1P U40 ( .A(Packet_In[5]), .Z(n127) );
  N1M1P U41 ( .A(Packet_In[10]), .Z(n137) );
  N1M1P U42 ( .A(Packet_In[25]), .Z(n151) );
  N1M1P U43 ( .A(Packet_In[6]), .Z(n129) );
  N1M1P U44 ( .A(Packet_In[4]), .Z(n125) );
  N1M1P U45 ( .A(Packet_In[14]), .Z(n145) );
  N1M1P U46 ( .A(Packet_In[11]), .Z(n139) );
  N1M1P U47 ( .A(Packet_In[7]), .Z(n131) );
  N1M1P U48 ( .A(Packet_In[9]), .Z(n135) );
  N1M1P U49 ( .A(Packet_In[12]), .Z(n141) );
  N1M1P U50 ( .A(Packet_In[26]), .Z(n153) );
  N1M1P U51 ( .A(Packet_In[15]), .Z(n147) );
  N1M1P U52 ( .A(Packet_In[24]), .Z(n149) );
  N1M1P U53 ( .A(Packet_In[1]), .Z(n119) );
  BUFM2P U54 ( .A(n162), .Z(n8) );
  N1M2P U55 ( .A(n7), .Z(n80) );
  OAI211M1P U56 ( .A(n113), .B(n112), .C(Rst_n), .D(n111), .Z(n163) );
  N1M2P U57 ( .A(n15), .Z(n112) );
  NR2M1P U58 ( .A(n110), .B(n7), .Z(n168) );
  NR2M1P U59 ( .A(n15), .B(n168), .Z(n167) );
  AOI22CDNM1P U60 ( .A(n167), .B(n20), .C(n167), .D(n20), .Z(n170) );
  N1M1P U61 ( .A(n168), .Z(n14) );
  AOI22M1P U62 ( .A(Count[0]), .B(n112), .C(n14), .D(n20), .Z(n11) );
  AOI22CDNM1P U63 ( .A(Count[1]), .B(n11), .C(n11), .D(Count[1]), .Z(n171) );
  ND3M1P U64 ( .A(n20), .B(n16), .C(n19), .Z(n49) );
  ND2M1P U65 ( .A(Count[1]), .B(Read_Ack), .Z(n10) );
  OAI211M1P U66 ( .A(Count[1]), .B(n112), .C(n11), .D(n10), .Z(n12) );
  AOI22M1P U67 ( .A(n15), .B(n113), .C(Count[2]), .D(n12), .Z(n13) );
  OAI21M1P U68 ( .A(n49), .B(n14), .C(n13), .Z(n172) );
  AOI22CDNM1P U69 ( .A(n17), .B(n166), .C(\Queue[4][31] ), .D(n17), .Z(n173)
         );
  AOI22CDNM1P U70 ( .A(n17), .B(n117), .C(\Queue[4][0] ), .D(n17), .Z(n174) );
  AOI22CDNM1P U71 ( .A(n17), .B(n119), .C(\Queue[4][1] ), .D(n17), .Z(n175) );
  AOI22CDNM1P U72 ( .A(n17), .B(n121), .C(\Queue[4][2] ), .D(n17), .Z(n176) );
  AOI22CDNM1P U73 ( .A(n17), .B(n123), .C(\Queue[4][3] ), .D(n17), .Z(n177) );
  AOI22CDNM1P U74 ( .A(n17), .B(n125), .C(\Queue[4][4] ), .D(n17), .Z(n178) );
  AOI22CDNM1P U75 ( .A(n17), .B(n127), .C(\Queue[4][5] ), .D(n17), .Z(n179) );
  AOI22CDNM1P U76 ( .A(n17), .B(n129), .C(\Queue[4][6] ), .D(n17), .Z(n180) );
  AOI22CDNM1P U77 ( .A(n17), .B(n131), .C(\Queue[4][7] ), .D(n17), .Z(n181) );
  AOI22CDNM1P U78 ( .A(n17), .B(n133), .C(\Queue[4][8] ), .D(n17), .Z(n182) );
  AOI22CDNM1P U79 ( .A(n17), .B(n135), .C(\Queue[4][9] ), .D(n17), .Z(n183) );
  AOI22CDNM1P U80 ( .A(n17), .B(n137), .C(\Queue[4][10] ), .D(n17), .Z(n184)
         );
  AOI22CDNM1P U81 ( .A(n17), .B(n139), .C(\Queue[4][11] ), .D(n17), .Z(n185)
         );
  AOI22CDNM1P U82 ( .A(n17), .B(n141), .C(\Queue[4][12] ), .D(n17), .Z(n186)
         );
  AOI22CDNM1P U83 ( .A(n17), .B(n143), .C(\Queue[4][13] ), .D(n17), .Z(n187)
         );
  AOI22CDNM1P U84 ( .A(n17), .B(n145), .C(\Queue[4][14] ), .D(n17), .Z(n188)
         );
  AOI22CDNM1P U85 ( .A(n17), .B(n147), .C(\Queue[4][15] ), .D(n17), .Z(n189)
         );
  AOI22CDNM1P U86 ( .A(n17), .B(n149), .C(\Queue[4][24] ), .D(n17), .Z(n190)
         );
  AOI22CDNM1P U87 ( .A(n17), .B(n151), .C(\Queue[4][25] ), .D(n17), .Z(n191)
         );
  AOI22CDNM1P U88 ( .A(n17), .B(n153), .C(\Queue[4][26] ), .D(n17), .Z(n192)
         );
  AOI22CDNM1P U89 ( .A(n17), .B(n155), .C(\Queue[4][27] ), .D(n17), .Z(n193)
         );
  AOI22CDNM1P U90 ( .A(n17), .B(n157), .C(\Queue[4][28] ), .D(n17), .Z(n194)
         );
  AOI22CDNM1P U91 ( .A(n17), .B(n159), .C(\Queue[4][29] ), .D(n17), .Z(n195)
         );
  AOI22CDNM1P U92 ( .A(n17), .B(n161), .C(\Queue[4][30] ), .D(n17), .Z(n196)
         );
  OAI22CDNM1P U93 ( .A(n112), .B(n18), .C(n167), .D(Full), .Z(n197) );
  OA21M1P U94 ( .A(n112), .B(n169), .C(Rst_n), .Z(n21) );
  AOI21M1P U95 ( .A(n7), .B(n81), .C(n114), .Z(n46) );
  AOI22M1P U96 ( .A(\Queue[2][0] ), .B(n6), .C(\Queue[1][0] ), .D(n3), .Z(n22)
         );
  OAI21M1P U97 ( .A(n117), .B(n48), .C(n22), .Z(n198) );
  AOI22M1P U98 ( .A(n6), .B(\Queue[2][1] ), .C(\Queue[1][1] ), .D(n3), .Z(n23)
         );
  OAI21M1P U99 ( .A(n48), .B(n119), .C(n23), .Z(n199) );
  AOI22M1P U100 ( .A(n6), .B(\Queue[2][2] ), .C(\Queue[1][2] ), .D(n3), .Z(n24) );
  OAI21M1P U101 ( .A(n48), .B(n121), .C(n24), .Z(n200) );
  AOI22M1P U102 ( .A(n6), .B(\Queue[2][3] ), .C(\Queue[1][3] ), .D(n3), .Z(n25) );
  OAI21M1P U103 ( .A(n48), .B(n123), .C(n25), .Z(n201) );
  AOI22M1P U104 ( .A(n6), .B(\Queue[2][4] ), .C(\Queue[1][4] ), .D(n3), .Z(n26) );
  OAI21M1P U105 ( .A(n48), .B(n125), .C(n26), .Z(n202) );
  AOI22M1P U106 ( .A(n6), .B(\Queue[2][5] ), .C(\Queue[1][5] ), .D(n3), .Z(n27) );
  OAI21M1P U107 ( .A(n48), .B(n127), .C(n27), .Z(n203) );
  AOI22M1P U108 ( .A(n6), .B(\Queue[2][6] ), .C(\Queue[1][6] ), .D(n3), .Z(n28) );
  OAI21M1P U109 ( .A(n48), .B(n129), .C(n28), .Z(n204) );
  AOI22M1P U110 ( .A(n6), .B(\Queue[2][7] ), .C(\Queue[1][7] ), .D(n3), .Z(n29) );
  OAI21M1P U111 ( .A(n48), .B(n131), .C(n29), .Z(n205) );
  AOI22M1P U112 ( .A(n6), .B(\Queue[2][8] ), .C(\Queue[1][8] ), .D(n3), .Z(n30) );
  OAI21M1P U113 ( .A(n48), .B(n133), .C(n30), .Z(n206) );
  AOI22M1P U114 ( .A(n6), .B(\Queue[2][9] ), .C(\Queue[1][9] ), .D(n45), .Z(
        n31) );
  OAI21M1P U115 ( .A(n48), .B(n135), .C(n31), .Z(n207) );
  AOI22M1P U116 ( .A(n6), .B(\Queue[2][10] ), .C(\Queue[1][10] ), .D(n45), .Z(
        n32) );
  OAI21M1P U117 ( .A(n48), .B(n137), .C(n32), .Z(n208) );
  AOI22M1P U118 ( .A(n6), .B(\Queue[2][11] ), .C(\Queue[1][11] ), .D(n45), .Z(
        n33) );
  OAI21M1P U119 ( .A(n48), .B(n139), .C(n33), .Z(n217) );
  AOI22M1P U120 ( .A(n6), .B(\Queue[2][12] ), .C(\Queue[1][12] ), .D(n45), .Z(
        n34) );
  OAI21M1P U121 ( .A(n48), .B(n141), .C(n34), .Z(n218) );
  AOI22M1P U122 ( .A(n6), .B(\Queue[2][13] ), .C(\Queue[1][13] ), .D(n45), .Z(
        n35) );
  OAI21M1P U123 ( .A(n48), .B(n143), .C(n35), .Z(n219) );
  AOI22M1P U124 ( .A(n6), .B(\Queue[2][14] ), .C(\Queue[1][14] ), .D(n45), .Z(
        n36) );
  OAI21M1P U125 ( .A(n48), .B(n145), .C(n36), .Z(n220) );
  AOI22M1P U126 ( .A(n6), .B(\Queue[2][15] ), .C(\Queue[1][15] ), .D(n45), .Z(
        n37) );
  OAI21M1P U127 ( .A(n48), .B(n147), .C(n37), .Z(n221) );
  AOI22M1P U128 ( .A(n6), .B(\Queue[2][24] ), .C(\Queue[1][24] ), .D(n3), .Z(
        n38) );
  OAI21M1P U129 ( .A(n48), .B(n149), .C(n38), .Z(n222) );
  AOI22M1P U130 ( .A(n6), .B(\Queue[2][25] ), .C(\Queue[1][25] ), .D(n3), .Z(
        n39) );
  OAI21M1P U131 ( .A(n48), .B(n151), .C(n39), .Z(n223) );
  AOI22M1P U132 ( .A(n6), .B(\Queue[2][26] ), .C(\Queue[1][26] ), .D(n3), .Z(
        n40) );
  OAI21M1P U133 ( .A(n48), .B(n153), .C(n40), .Z(n224) );
  AOI22M1P U134 ( .A(n6), .B(\Queue[2][27] ), .C(\Queue[1][27] ), .D(n3), .Z(
        n41) );
  OAI21M1P U135 ( .A(n48), .B(n155), .C(n41), .Z(n249) );
  AOI22M1P U136 ( .A(n6), .B(\Queue[2][28] ), .C(\Queue[1][28] ), .D(n3), .Z(
        n42) );
  OAI21M1P U137 ( .A(n48), .B(n157), .C(n42), .Z(n250) );
  AOI22M1P U138 ( .A(n6), .B(\Queue[2][29] ), .C(\Queue[1][29] ), .D(n3), .Z(
        n43) );
  OAI21M1P U139 ( .A(n48), .B(n159), .C(n43), .Z(n251) );
  AOI22M1P U140 ( .A(n6), .B(\Queue[2][30] ), .C(\Queue[1][30] ), .D(n3), .Z(
        n44) );
  OAI21M1P U141 ( .A(n48), .B(n161), .C(n44), .Z(n252) );
  AOI22M1P U142 ( .A(n6), .B(\Queue[2][31] ), .C(\Queue[1][31] ), .D(n3), .Z(
        n47) );
  OAI21M1P U143 ( .A(n48), .B(n166), .C(n47), .Z(n253) );
  OAI21M1P U144 ( .A(n50), .B(n49), .C(n114), .Z(n51) );
  AOI21M1P U145 ( .A(n7), .B(n169), .C(n114), .Z(n76) );
  AOI22M1P U146 ( .A(\Queue[1][0] ), .B(n4), .C(n75), .D(Packet_Out[0]), .Z(
        n52) );
  OAI21M1P U147 ( .A(n117), .B(n78), .C(n52), .Z(n254) );
  AOI22M1P U148 ( .A(\Queue[1][1] ), .B(n4), .C(n75), .D(Packet_Out[1]), .Z(
        n53) );
  OAI21M1P U149 ( .A(n119), .B(n78), .C(n53), .Z(n255) );
  AOI22M1P U150 ( .A(\Queue[1][2] ), .B(n4), .C(n75), .D(Packet_Out[2]), .Z(
        n54) );
  OAI21M1P U151 ( .A(n121), .B(n78), .C(n54), .Z(n256) );
  AOI22M1P U152 ( .A(\Queue[1][3] ), .B(n4), .C(n75), .D(Packet_Out[3]), .Z(
        n55) );
  OAI21M1P U153 ( .A(n123), .B(n78), .C(n55), .Z(n281) );
  AOI22M1P U154 ( .A(\Queue[1][4] ), .B(n4), .C(n75), .D(Packet_Out[4]), .Z(
        n56) );
  OAI21M1P U155 ( .A(n125), .B(n78), .C(n56), .Z(n282) );
  AOI22M1P U156 ( .A(\Queue[1][5] ), .B(n4), .C(n75), .D(Packet_Out[5]), .Z(
        n57) );
  OAI21M1P U157 ( .A(n127), .B(n78), .C(n57), .Z(n283) );
  AOI22M1P U158 ( .A(\Queue[1][6] ), .B(n4), .C(n75), .D(Packet_Out[6]), .Z(
        n58) );
  OAI21M1P U159 ( .A(n129), .B(n78), .C(n58), .Z(n284) );
  AOI22M1P U160 ( .A(\Queue[1][7] ), .B(n4), .C(n75), .D(Packet_Out[7]), .Z(
        n59) );
  OAI21M1P U161 ( .A(n131), .B(n78), .C(n59), .Z(n285) );
  AOI22M1P U162 ( .A(\Queue[1][8] ), .B(n4), .C(n75), .D(Packet_Out[8]), .Z(
        n60) );
  OAI21M1P U163 ( .A(n133), .B(n78), .C(n60), .Z(n286) );
  AOI22M1P U164 ( .A(\Queue[1][9] ), .B(n4), .C(n75), .D(Packet_Out[9]), .Z(
        n61) );
  OAI21M1P U165 ( .A(n135), .B(n78), .C(n61), .Z(n287) );
  AOI22M1P U166 ( .A(\Queue[1][10] ), .B(n4), .C(n75), .D(Packet_Out[10]), .Z(
        n62) );
  OAI21M1P U167 ( .A(n137), .B(n78), .C(n62), .Z(n288) );
  AOI22M1P U168 ( .A(\Queue[1][11] ), .B(n4), .C(n75), .D(Packet_Out[11]), .Z(
        n63) );
  OAI21M1P U169 ( .A(n139), .B(n78), .C(n63), .Z(n294) );
  AOI22M1P U170 ( .A(\Queue[1][12] ), .B(n4), .C(n75), .D(Packet_Out[12]), .Z(
        n64) );
  OAI21M1P U171 ( .A(n141), .B(n78), .C(n64), .Z(n295) );
  AOI22M1P U172 ( .A(\Queue[1][13] ), .B(n4), .C(n75), .D(Packet_Out[13]), .Z(
        n65) );
  OAI21M1P U173 ( .A(n143), .B(n78), .C(n65), .Z(n296) );
  AOI22M1P U174 ( .A(\Queue[1][14] ), .B(n4), .C(n75), .D(Packet_Out[14]), .Z(
        n66) );
  OAI21M1P U175 ( .A(n145), .B(n78), .C(n66), .Z(n297) );
  AOI22M1P U176 ( .A(\Queue[1][15] ), .B(n4), .C(n75), .D(Packet_Out[15]), .Z(
        n67) );
  OAI21M1P U177 ( .A(n147), .B(n78), .C(n67), .Z(n298) );
  AOI22M1P U178 ( .A(\Queue[1][24] ), .B(n4), .C(n75), .D(Packet_Out[24]), .Z(
        n68) );
  OAI21M1P U179 ( .A(n149), .B(n78), .C(n68), .Z(n299) );
  AOI22M1P U180 ( .A(\Queue[1][25] ), .B(n4), .C(n75), .D(Packet_Out[25]), .Z(
        n69) );
  OAI21M1P U181 ( .A(n151), .B(n78), .C(n69), .Z(n300) );
  AOI22M1P U182 ( .A(\Queue[1][26] ), .B(n4), .C(n75), .D(Packet_Out[26]), .Z(
        n70) );
  OAI21M1P U183 ( .A(n153), .B(n78), .C(n70), .Z(n301) );
  AOI22M1P U184 ( .A(\Queue[1][27] ), .B(n4), .C(n75), .D(Packet_Out[27]), .Z(
        n71) );
  OAI21M1P U185 ( .A(n155), .B(n78), .C(n71), .Z(n302) );
  AOI22M1P U186 ( .A(\Queue[1][28] ), .B(n4), .C(n75), .D(Packet_Out[28]), .Z(
        n72) );
  OAI21M1P U187 ( .A(n157), .B(n78), .C(n72), .Z(n303) );
  AOI22M1P U188 ( .A(\Queue[1][29] ), .B(n4), .C(n75), .D(Packet_Out[29]), .Z(
        n73) );
  OAI21M1P U189 ( .A(n159), .B(n78), .C(n73), .Z(n304) );
  AOI22M1P U190 ( .A(\Queue[1][30] ), .B(n4), .C(n75), .D(Packet_Out[30]), .Z(
        n74) );
  OAI21M1P U191 ( .A(n161), .B(n78), .C(n74), .Z(n305) );
  AOI22M1P U192 ( .A(\Queue[1][31] ), .B(n4), .C(n75), .D(Packet_Out[31]), .Z(
        n77) );
  OAI21M1P U193 ( .A(n166), .B(n78), .C(n77), .Z(n306) );
  OA21M1P U194 ( .A(n112), .B(n81), .C(Rst_n), .Z(n79) );
  ND2M1P U195 ( .A(n80), .B(n110), .Z(n111) );
  AOI21M1P U196 ( .A(n7), .B(n113), .C(n114), .Z(n105) );
  AOI22M1P U197 ( .A(\Queue[2][0] ), .B(n106), .C(\Queue[3][0] ), .D(n5), .Z(
        n82) );
  OAI21M1P U198 ( .A(n117), .B(n108), .C(n82), .Z(n307) );
  AOI22M1P U199 ( .A(\Queue[2][1] ), .B(n106), .C(n5), .D(\Queue[3][1] ), .Z(
        n83) );
  OAI21M1P U200 ( .A(n119), .B(n108), .C(n83), .Z(n308) );
  AOI22M1P U201 ( .A(\Queue[2][2] ), .B(n106), .C(n5), .D(\Queue[3][2] ), .Z(
        n84) );
  OAI21M1P U202 ( .A(n121), .B(n108), .C(n84), .Z(n309) );
  AOI22M1P U203 ( .A(\Queue[2][3] ), .B(n106), .C(n5), .D(\Queue[3][3] ), .Z(
        n85) );
  OAI21M1P U204 ( .A(n123), .B(n108), .C(n85), .Z(n310) );
  AOI22M1P U205 ( .A(\Queue[2][4] ), .B(n106), .C(n5), .D(\Queue[3][4] ), .Z(
        n86) );
  OAI21M1P U206 ( .A(n125), .B(n108), .C(n86), .Z(n311) );
  AOI22M1P U207 ( .A(\Queue[2][5] ), .B(n106), .C(n5), .D(\Queue[3][5] ), .Z(
        n87) );
  OAI21M1P U208 ( .A(n127), .B(n108), .C(n87), .Z(n312) );
  AOI22M1P U209 ( .A(\Queue[2][6] ), .B(n106), .C(n5), .D(\Queue[3][6] ), .Z(
        n88) );
  OAI21M1P U210 ( .A(n129), .B(n108), .C(n88), .Z(n313) );
  AOI22M1P U211 ( .A(\Queue[2][7] ), .B(n106), .C(n5), .D(\Queue[3][7] ), .Z(
        n89) );
  OAI21M1P U212 ( .A(n131), .B(n108), .C(n89), .Z(n314) );
  AOI22M1P U213 ( .A(\Queue[2][8] ), .B(n106), .C(n5), .D(\Queue[3][8] ), .Z(
        n90) );
  OAI21M1P U214 ( .A(n133), .B(n108), .C(n90), .Z(n315) );
  AOI22M1P U215 ( .A(\Queue[2][9] ), .B(n106), .C(n5), .D(\Queue[3][9] ), .Z(
        n91) );
  OAI21M1P U216 ( .A(n135), .B(n108), .C(n91), .Z(n316) );
  AOI22M1P U217 ( .A(\Queue[2][10] ), .B(n106), .C(n5), .D(\Queue[3][10] ), 
        .Z(n92) );
  OAI21M1P U218 ( .A(n137), .B(n108), .C(n92), .Z(n317) );
  AOI22M1P U219 ( .A(\Queue[2][11] ), .B(n106), .C(n5), .D(\Queue[3][11] ), 
        .Z(n93) );
  OAI21M1P U220 ( .A(n139), .B(n108), .C(n93), .Z(n318) );
  AOI22M1P U221 ( .A(\Queue[2][12] ), .B(n106), .C(n5), .D(\Queue[3][12] ), 
        .Z(n94) );
  OAI21M1P U222 ( .A(n141), .B(n108), .C(n94), .Z(n319) );
  AOI22M1P U223 ( .A(\Queue[2][13] ), .B(n106), .C(n5), .D(\Queue[3][13] ), 
        .Z(n95) );
  OAI21M1P U224 ( .A(n143), .B(n108), .C(n95), .Z(n320) );
  AOI22M1P U225 ( .A(\Queue[2][14] ), .B(n106), .C(n5), .D(\Queue[3][14] ), 
        .Z(n96) );
  OAI21M1P U226 ( .A(n145), .B(n108), .C(n96), .Z(n321) );
  AOI22M1P U227 ( .A(\Queue[2][15] ), .B(n106), .C(n5), .D(\Queue[3][15] ), 
        .Z(n97) );
  OAI21M1P U228 ( .A(n147), .B(n108), .C(n97), .Z(n322) );
  AOI22M1P U229 ( .A(\Queue[2][24] ), .B(n106), .C(n5), .D(\Queue[3][24] ), 
        .Z(n98) );
  OAI21M1P U230 ( .A(n149), .B(n108), .C(n98), .Z(n323) );
  AOI22M1P U231 ( .A(\Queue[2][25] ), .B(n106), .C(n5), .D(\Queue[3][25] ), 
        .Z(n99) );
  OAI21M1P U232 ( .A(n151), .B(n108), .C(n99), .Z(n324) );
  AOI22M1P U233 ( .A(\Queue[2][26] ), .B(n106), .C(n5), .D(\Queue[3][26] ), 
        .Z(n100) );
  OAI21M1P U234 ( .A(n153), .B(n108), .C(n100), .Z(n325) );
  AOI22M1P U235 ( .A(\Queue[2][27] ), .B(n106), .C(n5), .D(\Queue[3][27] ), 
        .Z(n101) );
  OAI21M1P U236 ( .A(n155), .B(n108), .C(n101), .Z(n326) );
  AOI22M1P U237 ( .A(\Queue[2][28] ), .B(n106), .C(n5), .D(\Queue[3][28] ), 
        .Z(n102) );
  OAI21M1P U238 ( .A(n157), .B(n108), .C(n102), .Z(n327) );
  AOI22M1P U239 ( .A(\Queue[2][29] ), .B(n106), .C(n5), .D(\Queue[3][29] ), 
        .Z(n103) );
  OAI21M1P U240 ( .A(n159), .B(n108), .C(n103), .Z(n328) );
  AOI22M1P U241 ( .A(\Queue[2][30] ), .B(n106), .C(n5), .D(\Queue[3][30] ), 
        .Z(n104) );
  OAI21M1P U242 ( .A(n161), .B(n108), .C(n104), .Z(n329) );
  AOI22M1P U243 ( .A(\Queue[2][31] ), .B(n106), .C(n5), .D(\Queue[3][31] ), 
        .Z(n107) );
  OAI21M1P U244 ( .A(n166), .B(n108), .C(n107), .Z(n330) );
  OA21M1P U245 ( .A(n112), .B(n113), .C(Rst_n), .Z(n109) );
  AOI22M1P U246 ( .A(\Queue[3][0] ), .B(n9), .C(n8), .D(\Queue[4][0] ), .Z(
        n116) );
  OAI21M1P U247 ( .A(n117), .B(n165), .C(n116), .Z(n331) );
  AOI22M1P U248 ( .A(\Queue[3][1] ), .B(n9), .C(n8), .D(\Queue[4][1] ), .Z(
        n118) );
  OAI21M1P U249 ( .A(n119), .B(n165), .C(n118), .Z(n332) );
  AOI22M1P U250 ( .A(\Queue[3][2] ), .B(n9), .C(n8), .D(\Queue[4][2] ), .Z(
        n120) );
  OAI21M1P U251 ( .A(n121), .B(n165), .C(n120), .Z(n333) );
  AOI22M1P U252 ( .A(\Queue[3][3] ), .B(n9), .C(n8), .D(\Queue[4][3] ), .Z(
        n122) );
  OAI21M1P U253 ( .A(n123), .B(n165), .C(n122), .Z(n334) );
  AOI22M1P U254 ( .A(\Queue[3][4] ), .B(n9), .C(n8), .D(\Queue[4][4] ), .Z(
        n124) );
  OAI21M1P U255 ( .A(n125), .B(n165), .C(n124), .Z(n335) );
  AOI22M1P U256 ( .A(\Queue[3][5] ), .B(n9), .C(n8), .D(\Queue[4][5] ), .Z(
        n126) );
  OAI21M1P U257 ( .A(n127), .B(n165), .C(n126), .Z(n336) );
  AOI22M1P U258 ( .A(\Queue[3][6] ), .B(n9), .C(n8), .D(\Queue[4][6] ), .Z(
        n128) );
  OAI21M1P U259 ( .A(n129), .B(n165), .C(n128), .Z(n337) );
  AOI22M1P U260 ( .A(\Queue[3][7] ), .B(n9), .C(n8), .D(\Queue[4][7] ), .Z(
        n130) );
  OAI21M1P U261 ( .A(n131), .B(n165), .C(n130), .Z(n338) );
  AOI22M1P U262 ( .A(\Queue[3][8] ), .B(n9), .C(n8), .D(\Queue[4][8] ), .Z(
        n132) );
  OAI21M1P U263 ( .A(n133), .B(n165), .C(n132), .Z(n339) );
  AOI22M1P U264 ( .A(\Queue[3][9] ), .B(n9), .C(n8), .D(\Queue[4][9] ), .Z(
        n134) );
  OAI21M1P U265 ( .A(n135), .B(n165), .C(n134), .Z(n340) );
  AOI22M1P U266 ( .A(\Queue[3][10] ), .B(n9), .C(n162), .D(\Queue[4][10] ), 
        .Z(n136) );
  OAI21M1P U267 ( .A(n137), .B(n165), .C(n136), .Z(n341) );
  AOI22M1P U268 ( .A(\Queue[3][11] ), .B(n9), .C(n162), .D(\Queue[4][11] ), 
        .Z(n138) );
  OAI21M1P U269 ( .A(n139), .B(n165), .C(n138), .Z(n342) );
  AOI22M1P U270 ( .A(\Queue[3][12] ), .B(n9), .C(n162), .D(\Queue[4][12] ), 
        .Z(n140) );
  OAI21M1P U271 ( .A(n141), .B(n165), .C(n140), .Z(n343) );
  AOI22M1P U272 ( .A(\Queue[3][13] ), .B(n9), .C(n162), .D(\Queue[4][13] ), 
        .Z(n142) );
  OAI21M1P U273 ( .A(n143), .B(n165), .C(n142), .Z(n344) );
  AOI22M1P U274 ( .A(\Queue[3][14] ), .B(n9), .C(n162), .D(\Queue[4][14] ), 
        .Z(n144) );
  OAI21M1P U275 ( .A(n145), .B(n165), .C(n144), .Z(n345) );
  AOI22M1P U276 ( .A(\Queue[3][15] ), .B(n9), .C(n162), .D(\Queue[4][15] ), 
        .Z(n146) );
  OAI21M1P U277 ( .A(n147), .B(n165), .C(n146), .Z(n346) );
  AOI22M1P U278 ( .A(\Queue[3][24] ), .B(n9), .C(n162), .D(\Queue[4][24] ), 
        .Z(n148) );
  OAI21M1P U279 ( .A(n149), .B(n165), .C(n148), .Z(n347) );
  AOI22M1P U280 ( .A(\Queue[3][25] ), .B(n9), .C(n162), .D(\Queue[4][25] ), 
        .Z(n150) );
  OAI21M1P U281 ( .A(n151), .B(n165), .C(n150), .Z(n348) );
  AOI22M1P U282 ( .A(\Queue[3][26] ), .B(n9), .C(n162), .D(\Queue[4][26] ), 
        .Z(n152) );
  OAI21M1P U283 ( .A(n153), .B(n165), .C(n152), .Z(n349) );
  AOI22M1P U284 ( .A(\Queue[3][27] ), .B(n9), .C(n162), .D(\Queue[4][27] ), 
        .Z(n154) );
  OAI21M1P U285 ( .A(n155), .B(n165), .C(n154), .Z(n350) );
  AOI22M1P U286 ( .A(\Queue[3][28] ), .B(n163), .C(n162), .D(\Queue[4][28] ), 
        .Z(n156) );
  OAI21M1P U287 ( .A(n157), .B(n165), .C(n156), .Z(n351) );
  AOI22M1P U288 ( .A(\Queue[3][29] ), .B(n163), .C(n162), .D(\Queue[4][29] ), 
        .Z(n158) );
  OAI21M1P U289 ( .A(n159), .B(n165), .C(n158), .Z(n352) );
  AOI22M1P U290 ( .A(\Queue[3][30] ), .B(n163), .C(n8), .D(\Queue[4][30] ), 
        .Z(n160) );
  OAI21M1P U291 ( .A(n161), .B(n165), .C(n160), .Z(n353) );
  AOI22M1P U292 ( .A(\Queue[3][31] ), .B(n9), .C(n8), .D(\Queue[4][31] ), .Z(
        n164) );
  OAI21M1P U293 ( .A(n166), .B(n165), .C(n164), .Z(n354) );
  N1M1P U294 ( .A(n355), .Z(Empty) );
  AOI22M1P U295 ( .A(n169), .B(n168), .C(n167), .D(Empty), .Z(n356) );
endmodule


module Node_Manager ( Clk_r, Rst_n, Packet_From_Core, Packet_From_Node, 
        Packet_From_Node_Valid, Read_Packet, To_Node_Write, Router_Address, 
        Link_Config, Packet_To_Core, Packet_To_Node, Packet_To_Node_Valid, 
        Core_Load_Ack, Queue_Empty, To_Node_Full );
  input [31:0] Packet_From_Core;
  input [31:0] Packet_From_Node;
  output [7:0] Router_Address;
  output [3:0] Link_Config;
  output [31:0] Packet_To_Core;
  output [31:0] Packet_To_Node;
  input Clk_r, Rst_n, Packet_From_Node_Valid, Read_Packet, To_Node_Write;
  output Packet_To_Node_Valid, Core_Load_Ack, Queue_Empty, To_Node_Full;
  wire   Write_Queue, Queue_Full, Read_Out_Queue, Out_Queue_Empty, N8, N42,
         N43, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7;

  Packet_Queue_2 In_Queue ( .Clk_r(Clk_r), .Rst_n(Rst_n), .Packet_In({
        Packet_From_Node[31:24], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, Packet_From_Node[15:0]}), .Read_Ack(Read_Packet), .Write_Ack(
        Write_Queue), .Packet_Out({Packet_To_Core[31:24], 
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, Packet_To_Core[15:0]}), .Empty(Queue_Empty), .Full(Queue_Full) );
  Packet_Queue_1 Out_Queue ( .Clk_r(Clk_r), .Rst_n(Rst_n), .Packet_In(
        Packet_From_Core), .Read_Ack(Read_Out_Queue), .Write_Ack(To_Node_Write), .Packet_Out(Packet_To_Node), .Empty(Out_Queue_Empty), .Full(To_Node_Full) );
  FD2LQM1P \Router_Address_reg[0]  ( .D(Packet_From_Node[0]), .LD(n2), .CP(
        Clk_r), .CD(Rst_n), .Q(Router_Address[0]) );
  FD2LQM1P \Router_Address_reg[1]  ( .D(Packet_From_Node[1]), .LD(n2), .CP(
        Clk_r), .CD(Rst_n), .Q(Router_Address[1]) );
  FD2LQM1P \Router_Address_reg[2]  ( .D(Packet_From_Node[2]), .LD(n2), .CP(
        Clk_r), .CD(Rst_n), .Q(Router_Address[2]) );
  FD2LQM1P \Router_Address_reg[3]  ( .D(Packet_From_Node[3]), .LD(n2), .CP(
        Clk_r), .CD(Rst_n), .Q(Router_Address[3]) );
  FD2LQM1P \Router_Address_reg[4]  ( .D(Packet_From_Node[4]), .LD(n2), .CP(
        Clk_r), .CD(Rst_n), .Q(Router_Address[4]) );
  FD2LQM1P \Router_Address_reg[5]  ( .D(Packet_From_Node[5]), .LD(n2), .CP(
        Clk_r), .CD(Rst_n), .Q(Router_Address[5]) );
  FD2LQM1P \Router_Address_reg[6]  ( .D(Packet_From_Node[6]), .LD(n2), .CP(
        Clk_r), .CD(Rst_n), .Q(Router_Address[6]) );
  FD2LQM1P \Router_Address_reg[7]  ( .D(Packet_From_Node[7]), .LD(n2), .CP(
        Clk_r), .CD(Rst_n), .Q(Router_Address[7]) );
  FD2LQM1P \Link_Config_reg[0]  ( .D(Packet_From_Node[0]), .LD(n1), .CP(Clk_r), 
        .CD(Rst_n), .Q(Link_Config[0]) );
  FD2LQM1P \Link_Config_reg[1]  ( .D(Packet_From_Node[1]), .LD(n1), .CP(Clk_r), 
        .CD(Rst_n), .Q(Link_Config[1]) );
  FD2LQM1P \Link_Config_reg[2]  ( .D(Packet_From_Node[2]), .LD(n1), .CP(Clk_r), 
        .CD(Rst_n), .Q(Link_Config[2]) );
  FD2LQM1P \Link_Config_reg[3]  ( .D(Packet_From_Node[3]), .LD(n1), .CP(Clk_r), 
        .CD(Rst_n), .Q(Link_Config[3]) );
  FD2QM1P Read_Out_Queue_reg ( .D(Packet_To_Node_Valid), .CP(Clk_r), .CD(Rst_n), .Q(Read_Out_Queue) );
  FD2QM1P Packet_To_Node_Valid_reg ( .D(N8), .CP(Clk_r), .CD(Rst_n), .Q(
        Packet_To_Node_Valid) );
  FD2QM1P Core_Load_Ack_reg ( .D(N42), .CP(Clk_r), .CD(Rst_n), .Q(
        Core_Load_Ack) );
  FD2QM1P Write_Queue_reg ( .D(N43), .CP(Clk_r), .CD(Rst_n), .Q(Write_Queue)
         );
  NR2M1P U3 ( .A(Packet_From_Node[16]), .B(n10), .Z(n2) );
  ND4M1P U5 ( .A(Packet_From_Node[30]), .B(Packet_From_Node[31]), .C(
        Packet_From_Node[28]), .D(Packet_From_Node[29]), .Z(n5) );
  ND4M1P U6 ( .A(Packet_From_Node[26]), .B(Packet_From_Node[27]), .C(
        Packet_From_Node[24]), .D(Packet_From_Node[25]), .Z(n4) );
  AND2M1P U7 ( .A(n5), .B(n4), .Z(n3) );
  ND2BNM1P U8 ( .B(Core_Load_Ack), .A(Packet_From_Node_Valid), .Z(n6) );
  AOI21M1P U9 ( .A(n3), .B(Queue_Full), .C(n6), .Z(N42) );
  NR3CNM1P U10 ( .C(n3), .A(Queue_Full), .B(n6), .Z(N43) );
  NR2M1P U11 ( .A(Out_Queue_Empty), .B(Packet_To_Node_Valid), .Z(N8) );
  NR3M1P U12 ( .A(Packet_From_Node[23]), .B(Packet_From_Node[18]), .C(
        Packet_From_Node[17]), .Z(n9) );
  NR3M1P U13 ( .A(Packet_From_Node[19]), .B(Packet_From_Node[20]), .C(n4), .Z(
        n8) );
  NR3M1P U14 ( .A(Packet_From_Node[21]), .B(n6), .C(n5), .Z(n7) );
  ND4DNM1P U15 ( .D(Packet_From_Node[22]), .A(n9), .B(n8), .C(n7), .Z(n10) );
  NR2BNM1P U16 ( .B(Packet_From_Node[16]), .A(n10), .Z(n1) );
endmodule


module Packet_Queue_3 ( Clk_r, Rst_n, Packet_In, Read_Ack, Write_Ack, 
        Packet_Out, Empty, Full );
  input [31:0] Packet_In;
  output [31:0] Packet_Out;
  input Clk_r, Rst_n, Read_Ack, Write_Ack;
  output Empty, Full;
  wire   \Queue[4][31] , \Queue[4][30] , \Queue[4][29] , \Queue[4][28] ,
         \Queue[4][27] , \Queue[4][26] , \Queue[4][25] , \Queue[4][24] ,
         \Queue[4][23] , \Queue[4][22] , \Queue[4][21] , \Queue[4][20] ,
         \Queue[4][19] , \Queue[4][18] , \Queue[4][17] , \Queue[4][16] ,
         \Queue[4][15] , \Queue[4][14] , \Queue[4][13] , \Queue[4][12] ,
         \Queue[4][11] , \Queue[4][10] , \Queue[4][9] , \Queue[4][8] ,
         \Queue[4][7] , \Queue[4][6] , \Queue[4][5] , \Queue[4][4] ,
         \Queue[4][3] , \Queue[4][2] , \Queue[4][1] , \Queue[4][0] ,
         \Queue[3][31] , \Queue[3][30] , \Queue[3][29] , \Queue[3][28] ,
         \Queue[3][27] , \Queue[3][26] , \Queue[3][25] , \Queue[3][24] ,
         \Queue[3][23] , \Queue[3][22] , \Queue[3][21] , \Queue[3][20] ,
         \Queue[3][19] , \Queue[3][18] , \Queue[3][17] , \Queue[3][16] ,
         \Queue[3][15] , \Queue[3][14] , \Queue[3][13] , \Queue[3][12] ,
         \Queue[3][11] , \Queue[3][10] , \Queue[3][9] , \Queue[3][8] ,
         \Queue[3][7] , \Queue[3][6] , \Queue[3][5] , \Queue[3][4] ,
         \Queue[3][3] , \Queue[3][2] , \Queue[3][1] , \Queue[3][0] ,
         \Queue[2][31] , \Queue[2][30] , \Queue[2][29] , \Queue[2][28] ,
         \Queue[2][27] , \Queue[2][26] , \Queue[2][25] , \Queue[2][24] ,
         \Queue[2][23] , \Queue[2][22] , \Queue[2][21] , \Queue[2][20] ,
         \Queue[2][19] , \Queue[2][18] , \Queue[2][17] , \Queue[2][16] ,
         \Queue[2][15] , \Queue[2][14] , \Queue[2][13] , \Queue[2][12] ,
         \Queue[2][11] , \Queue[2][10] , \Queue[2][9] , \Queue[2][8] ,
         \Queue[2][7] , \Queue[2][6] , \Queue[2][5] , \Queue[2][4] ,
         \Queue[2][3] , \Queue[2][2] , \Queue[2][1] , \Queue[2][0] ,
         \Queue[1][31] , \Queue[1][30] , \Queue[1][29] , \Queue[1][28] ,
         \Queue[1][27] , \Queue[1][26] , \Queue[1][25] , \Queue[1][24] ,
         \Queue[1][23] , \Queue[1][22] , \Queue[1][21] , \Queue[1][20] ,
         \Queue[1][19] , \Queue[1][18] , \Queue[1][17] , \Queue[1][16] ,
         \Queue[1][15] , \Queue[1][14] , \Queue[1][13] , \Queue[1][12] ,
         \Queue[1][11] , \Queue[1][10] , \Queue[1][9] , \Queue[1][8] ,
         \Queue[1][7] , \Queue[1][6] , \Queue[1][5] , \Queue[1][4] ,
         \Queue[1][3] , \Queue[1][2] , \Queue[1][1] , \Queue[1][0] , n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542;
  wire   [2:0] Count;

  FDN2QM1P \Count_reg[0]  ( .D(n377), .CPN(Clk_r), .CD(Rst_n), .Q(Count[0]) );
  FDN2QM1P \Count_reg[1]  ( .D(n378), .CPN(Clk_r), .CD(Rst_n), .Q(Count[1]) );
  FDN2QM1P \Count_reg[2]  ( .D(n379), .CPN(Clk_r), .CD(Rst_n), .Q(Count[2]) );
  FDN1QM1P \Queue_reg[4][30]  ( .D(n411), .CPN(Clk_r), .Q(\Queue[4][30] ) );
  FDN1QM1P \Queue_reg[3][30]  ( .D(n539), .CPN(Clk_r), .Q(\Queue[3][30] ) );
  FDN1QM1P \Queue_reg[2][30]  ( .D(n507), .CPN(Clk_r), .Q(\Queue[2][30] ) );
  FDN1QM1P \Queue_reg[4][29]  ( .D(n410), .CPN(Clk_r), .Q(\Queue[4][29] ) );
  FDN1QM1P \Queue_reg[3][29]  ( .D(n538), .CPN(Clk_r), .Q(\Queue[3][29] ) );
  FDN1QM1P \Queue_reg[2][29]  ( .D(n506), .CPN(Clk_r), .Q(\Queue[2][29] ) );
  FDN1QM1P \Queue_reg[4][28]  ( .D(n409), .CPN(Clk_r), .Q(\Queue[4][28] ) );
  FDN1QM1P \Queue_reg[3][28]  ( .D(n537), .CPN(Clk_r), .Q(\Queue[3][28] ) );
  FDN1QM1P \Queue_reg[2][28]  ( .D(n505), .CPN(Clk_r), .Q(\Queue[2][28] ) );
  FDN1QM1P \Queue_reg[4][27]  ( .D(n408), .CPN(Clk_r), .Q(\Queue[4][27] ) );
  FDN1QM1P \Queue_reg[3][27]  ( .D(n536), .CPN(Clk_r), .Q(\Queue[3][27] ) );
  FDN1QM1P \Queue_reg[2][27]  ( .D(n504), .CPN(Clk_r), .Q(\Queue[2][27] ) );
  FDN1QM1P \Queue_reg[4][26]  ( .D(n407), .CPN(Clk_r), .Q(\Queue[4][26] ) );
  FDN1QM1P \Queue_reg[3][26]  ( .D(n535), .CPN(Clk_r), .Q(\Queue[3][26] ) );
  FDN1QM1P \Queue_reg[2][26]  ( .D(n503), .CPN(Clk_r), .Q(\Queue[2][26] ) );
  FDN1QM1P \Queue_reg[4][25]  ( .D(n406), .CPN(Clk_r), .Q(\Queue[4][25] ) );
  FDN1QM1P \Queue_reg[3][25]  ( .D(n534), .CPN(Clk_r), .Q(\Queue[3][25] ) );
  FDN1QM1P \Queue_reg[2][25]  ( .D(n502), .CPN(Clk_r), .Q(\Queue[2][25] ) );
  FDN1QM1P \Queue_reg[4][24]  ( .D(n405), .CPN(Clk_r), .Q(\Queue[4][24] ) );
  FDN1QM1P \Queue_reg[3][24]  ( .D(n533), .CPN(Clk_r), .Q(\Queue[3][24] ) );
  FDN1QM1P \Queue_reg[2][24]  ( .D(n501), .CPN(Clk_r), .Q(\Queue[2][24] ) );
  FDN1QM1P \Queue_reg[4][23]  ( .D(n404), .CPN(Clk_r), .Q(\Queue[4][23] ) );
  FDN1QM1P \Queue_reg[3][23]  ( .D(n532), .CPN(Clk_r), .Q(\Queue[3][23] ) );
  FDN1QM1P \Queue_reg[2][23]  ( .D(n500), .CPN(Clk_r), .Q(\Queue[2][23] ) );
  FDN1QM1P \Queue_reg[4][22]  ( .D(n403), .CPN(Clk_r), .Q(\Queue[4][22] ) );
  FDN1QM1P \Queue_reg[3][22]  ( .D(n531), .CPN(Clk_r), .Q(\Queue[3][22] ) );
  FDN1QM1P \Queue_reg[2][22]  ( .D(n499), .CPN(Clk_r), .Q(\Queue[2][22] ) );
  FDN1QM1P \Queue_reg[4][21]  ( .D(n402), .CPN(Clk_r), .Q(\Queue[4][21] ) );
  FDN1QM1P \Queue_reg[3][21]  ( .D(n530), .CPN(Clk_r), .Q(\Queue[3][21] ) );
  FDN1QM1P \Queue_reg[2][21]  ( .D(n498), .CPN(Clk_r), .Q(\Queue[2][21] ) );
  FDN1QM1P \Queue_reg[4][20]  ( .D(n401), .CPN(Clk_r), .Q(\Queue[4][20] ) );
  FDN1QM1P \Queue_reg[3][20]  ( .D(n529), .CPN(Clk_r), .Q(\Queue[3][20] ) );
  FDN1QM1P \Queue_reg[2][20]  ( .D(n497), .CPN(Clk_r), .Q(\Queue[2][20] ) );
  FDN1QM1P \Queue_reg[4][19]  ( .D(n400), .CPN(Clk_r), .Q(\Queue[4][19] ) );
  FDN1QM1P \Queue_reg[3][19]  ( .D(n528), .CPN(Clk_r), .Q(\Queue[3][19] ) );
  FDN1QM1P \Queue_reg[2][19]  ( .D(n496), .CPN(Clk_r), .Q(\Queue[2][19] ) );
  FDN1QM1P \Queue_reg[4][18]  ( .D(n399), .CPN(Clk_r), .Q(\Queue[4][18] ) );
  FDN1QM1P \Queue_reg[3][18]  ( .D(n527), .CPN(Clk_r), .Q(\Queue[3][18] ) );
  FDN1QM1P \Queue_reg[2][18]  ( .D(n495), .CPN(Clk_r), .Q(\Queue[2][18] ) );
  FDN1QM1P \Queue_reg[4][17]  ( .D(n398), .CPN(Clk_r), .Q(\Queue[4][17] ) );
  FDN1QM1P \Queue_reg[3][17]  ( .D(n526), .CPN(Clk_r), .Q(\Queue[3][17] ) );
  FDN1QM1P \Queue_reg[2][17]  ( .D(n494), .CPN(Clk_r), .Q(\Queue[2][17] ) );
  FDN1QM1P \Queue_reg[4][16]  ( .D(n397), .CPN(Clk_r), .Q(\Queue[4][16] ) );
  FDN1QM1P \Queue_reg[3][16]  ( .D(n525), .CPN(Clk_r), .Q(\Queue[3][16] ) );
  FDN1QM1P \Queue_reg[2][16]  ( .D(n493), .CPN(Clk_r), .Q(\Queue[2][16] ) );
  FDN1QM1P \Queue_reg[4][15]  ( .D(n396), .CPN(Clk_r), .Q(\Queue[4][15] ) );
  FDN1QM1P \Queue_reg[3][15]  ( .D(n524), .CPN(Clk_r), .Q(\Queue[3][15] ) );
  FDN1QM1P \Queue_reg[2][15]  ( .D(n492), .CPN(Clk_r), .Q(\Queue[2][15] ) );
  FDN1QM1P \Queue_reg[4][14]  ( .D(n395), .CPN(Clk_r), .Q(\Queue[4][14] ) );
  FDN1QM1P \Queue_reg[3][14]  ( .D(n523), .CPN(Clk_r), .Q(\Queue[3][14] ) );
  FDN1QM1P \Queue_reg[2][14]  ( .D(n491), .CPN(Clk_r), .Q(\Queue[2][14] ) );
  FDN1QM1P \Queue_reg[4][13]  ( .D(n394), .CPN(Clk_r), .Q(\Queue[4][13] ) );
  FDN1QM1P \Queue_reg[3][13]  ( .D(n522), .CPN(Clk_r), .Q(\Queue[3][13] ) );
  FDN1QM1P \Queue_reg[2][13]  ( .D(n490), .CPN(Clk_r), .Q(\Queue[2][13] ) );
  FDN1QM1P \Queue_reg[4][12]  ( .D(n393), .CPN(Clk_r), .Q(\Queue[4][12] ) );
  FDN1QM1P \Queue_reg[3][12]  ( .D(n521), .CPN(Clk_r), .Q(\Queue[3][12] ) );
  FDN1QM1P \Queue_reg[2][12]  ( .D(n489), .CPN(Clk_r), .Q(\Queue[2][12] ) );
  FDN1QM1P \Queue_reg[4][11]  ( .D(n392), .CPN(Clk_r), .Q(\Queue[4][11] ) );
  FDN1QM1P \Queue_reg[3][11]  ( .D(n520), .CPN(Clk_r), .Q(\Queue[3][11] ) );
  FDN1QM1P \Queue_reg[2][11]  ( .D(n488), .CPN(Clk_r), .Q(\Queue[2][11] ) );
  FDN1QM1P \Queue_reg[4][10]  ( .D(n391), .CPN(Clk_r), .Q(\Queue[4][10] ) );
  FDN1QM1P \Queue_reg[3][10]  ( .D(n519), .CPN(Clk_r), .Q(\Queue[3][10] ) );
  FDN1QM1P \Queue_reg[2][10]  ( .D(n487), .CPN(Clk_r), .Q(\Queue[2][10] ) );
  FDN1QM1P \Queue_reg[4][9]  ( .D(n390), .CPN(Clk_r), .Q(\Queue[4][9] ) );
  FDN1QM1P \Queue_reg[3][9]  ( .D(n518), .CPN(Clk_r), .Q(\Queue[3][9] ) );
  FDN1QM1P \Queue_reg[2][9]  ( .D(n486), .CPN(Clk_r), .Q(\Queue[2][9] ) );
  FDN1QM1P \Queue_reg[4][8]  ( .D(n389), .CPN(Clk_r), .Q(\Queue[4][8] ) );
  FDN1QM1P \Queue_reg[3][8]  ( .D(n517), .CPN(Clk_r), .Q(\Queue[3][8] ) );
  FDN1QM1P \Queue_reg[2][8]  ( .D(n485), .CPN(Clk_r), .Q(\Queue[2][8] ) );
  FDN1QM1P \Queue_reg[4][7]  ( .D(n388), .CPN(Clk_r), .Q(\Queue[4][7] ) );
  FDN1QM1P \Queue_reg[3][7]  ( .D(n516), .CPN(Clk_r), .Q(\Queue[3][7] ) );
  FDN1QM1P \Queue_reg[2][7]  ( .D(n484), .CPN(Clk_r), .Q(\Queue[2][7] ) );
  FDN1QM1P \Queue_reg[4][6]  ( .D(n387), .CPN(Clk_r), .Q(\Queue[4][6] ) );
  FDN1QM1P \Queue_reg[3][6]  ( .D(n515), .CPN(Clk_r), .Q(\Queue[3][6] ) );
  FDN1QM1P \Queue_reg[2][6]  ( .D(n483), .CPN(Clk_r), .Q(\Queue[2][6] ) );
  FDN1QM1P \Queue_reg[4][5]  ( .D(n386), .CPN(Clk_r), .Q(\Queue[4][5] ) );
  FDN1QM1P \Queue_reg[3][5]  ( .D(n514), .CPN(Clk_r), .Q(\Queue[3][5] ) );
  FDN1QM1P \Queue_reg[2][5]  ( .D(n482), .CPN(Clk_r), .Q(\Queue[2][5] ) );
  FDN1QM1P \Queue_reg[4][4]  ( .D(n385), .CPN(Clk_r), .Q(\Queue[4][4] ) );
  FDN1QM1P \Queue_reg[3][4]  ( .D(n513), .CPN(Clk_r), .Q(\Queue[3][4] ) );
  FDN1QM1P \Queue_reg[2][4]  ( .D(n481), .CPN(Clk_r), .Q(\Queue[2][4] ) );
  FDN1QM1P \Queue_reg[4][3]  ( .D(n384), .CPN(Clk_r), .Q(\Queue[4][3] ) );
  FDN1QM1P \Queue_reg[3][3]  ( .D(n512), .CPN(Clk_r), .Q(\Queue[3][3] ) );
  FDN1QM1P \Queue_reg[2][3]  ( .D(n480), .CPN(Clk_r), .Q(\Queue[2][3] ) );
  FDN1QM1P \Queue_reg[4][2]  ( .D(n383), .CPN(Clk_r), .Q(\Queue[4][2] ) );
  FDN1QM1P \Queue_reg[3][2]  ( .D(n511), .CPN(Clk_r), .Q(\Queue[3][2] ) );
  FDN1QM1P \Queue_reg[2][2]  ( .D(n479), .CPN(Clk_r), .Q(\Queue[2][2] ) );
  FDN1QM1P \Queue_reg[4][1]  ( .D(n382), .CPN(Clk_r), .Q(\Queue[4][1] ) );
  FDN1QM1P \Queue_reg[3][1]  ( .D(n510), .CPN(Clk_r), .Q(\Queue[3][1] ) );
  FDN1QM1P \Queue_reg[2][1]  ( .D(n478), .CPN(Clk_r), .Q(\Queue[2][1] ) );
  FDN1QM1P \Queue_reg[4][0]  ( .D(n381), .CPN(Clk_r), .Q(\Queue[4][0] ) );
  FDN1QM1P \Queue_reg[3][0]  ( .D(n509), .CPN(Clk_r), .Q(\Queue[3][0] ) );
  FDN1QM1P \Queue_reg[2][0]  ( .D(n477), .CPN(Clk_r), .Q(\Queue[2][0] ) );
  FDN1QM1P \Queue_reg[4][31]  ( .D(n380), .CPN(Clk_r), .Q(\Queue[4][31] ) );
  FDN1QM1P \Queue_reg[3][31]  ( .D(n540), .CPN(Clk_r), .Q(\Queue[3][31] ) );
  FDN1QM1P \Queue_reg[2][31]  ( .D(n508), .CPN(Clk_r), .Q(\Queue[2][31] ) );
  FDN2QM1P Full_reg ( .D(n412), .CPN(Clk_r), .CD(Rst_n), .Q(Full) );
  FDN1QM1P \Queue_reg[1][31]  ( .D(n444), .CPN(Clk_r), .Q(\Queue[1][31] ) );
  FDN1QM1P \Queue_reg[0][31]  ( .D(n476), .CPN(Clk_r), .Q(Packet_Out[31]) );
  FDN1QM1P \Queue_reg[1][30]  ( .D(n443), .CPN(Clk_r), .Q(\Queue[1][30] ) );
  FDN1QM1P \Queue_reg[0][30]  ( .D(n475), .CPN(Clk_r), .Q(Packet_Out[30]) );
  FDN1QM1P \Queue_reg[1][29]  ( .D(n442), .CPN(Clk_r), .Q(\Queue[1][29] ) );
  FDN1QM1P \Queue_reg[0][29]  ( .D(n474), .CPN(Clk_r), .Q(Packet_Out[29]) );
  FDN1QM1P \Queue_reg[1][28]  ( .D(n441), .CPN(Clk_r), .Q(\Queue[1][28] ) );
  FDN1QM1P \Queue_reg[0][28]  ( .D(n473), .CPN(Clk_r), .Q(Packet_Out[28]) );
  FDN1QM1P \Queue_reg[1][27]  ( .D(n440), .CPN(Clk_r), .Q(\Queue[1][27] ) );
  FDN1QM1P \Queue_reg[0][27]  ( .D(n472), .CPN(Clk_r), .Q(Packet_Out[27]) );
  FDN1QM1P \Queue_reg[1][26]  ( .D(n439), .CPN(Clk_r), .Q(\Queue[1][26] ) );
  FDN1QM1P \Queue_reg[0][26]  ( .D(n471), .CPN(Clk_r), .Q(Packet_Out[26]) );
  FDN1QM1P \Queue_reg[1][25]  ( .D(n438), .CPN(Clk_r), .Q(\Queue[1][25] ) );
  FDN1QM1P \Queue_reg[0][25]  ( .D(n470), .CPN(Clk_r), .Q(Packet_Out[25]) );
  FDN1QM1P \Queue_reg[1][24]  ( .D(n437), .CPN(Clk_r), .Q(\Queue[1][24] ) );
  FDN1QM1P \Queue_reg[0][24]  ( .D(n469), .CPN(Clk_r), .Q(Packet_Out[24]) );
  FDN1QM1P \Queue_reg[1][23]  ( .D(n436), .CPN(Clk_r), .Q(\Queue[1][23] ) );
  FDN1QM1P \Queue_reg[0][23]  ( .D(n468), .CPN(Clk_r), .Q(Packet_Out[23]) );
  FDN1QM1P \Queue_reg[1][22]  ( .D(n435), .CPN(Clk_r), .Q(\Queue[1][22] ) );
  FDN1QM1P \Queue_reg[0][22]  ( .D(n467), .CPN(Clk_r), .Q(Packet_Out[22]) );
  FDN1QM1P \Queue_reg[1][21]  ( .D(n434), .CPN(Clk_r), .Q(\Queue[1][21] ) );
  FDN1QM1P \Queue_reg[0][21]  ( .D(n466), .CPN(Clk_r), .Q(Packet_Out[21]) );
  FDN1QM1P \Queue_reg[1][20]  ( .D(n433), .CPN(Clk_r), .Q(\Queue[1][20] ) );
  FDN1QM1P \Queue_reg[0][20]  ( .D(n465), .CPN(Clk_r), .Q(Packet_Out[20]) );
  FDN1QM1P \Queue_reg[1][19]  ( .D(n432), .CPN(Clk_r), .Q(\Queue[1][19] ) );
  FDN1QM1P \Queue_reg[0][19]  ( .D(n464), .CPN(Clk_r), .Q(Packet_Out[19]) );
  FDN1QM1P \Queue_reg[1][18]  ( .D(n431), .CPN(Clk_r), .Q(\Queue[1][18] ) );
  FDN1QM1P \Queue_reg[0][18]  ( .D(n463), .CPN(Clk_r), .Q(Packet_Out[18]) );
  FDN1QM1P \Queue_reg[1][17]  ( .D(n430), .CPN(Clk_r), .Q(\Queue[1][17] ) );
  FDN1QM1P \Queue_reg[0][17]  ( .D(n462), .CPN(Clk_r), .Q(Packet_Out[17]) );
  FDN1QM1P \Queue_reg[1][16]  ( .D(n429), .CPN(Clk_r), .Q(\Queue[1][16] ) );
  FDN1QM1P \Queue_reg[0][16]  ( .D(n461), .CPN(Clk_r), .Q(Packet_Out[16]) );
  FDN1QM1P \Queue_reg[1][15]  ( .D(n428), .CPN(Clk_r), .Q(\Queue[1][15] ) );
  FDN1QM1P \Queue_reg[0][15]  ( .D(n460), .CPN(Clk_r), .Q(Packet_Out[15]) );
  FDN1QM1P \Queue_reg[1][14]  ( .D(n427), .CPN(Clk_r), .Q(\Queue[1][14] ) );
  FDN1QM1P \Queue_reg[0][14]  ( .D(n459), .CPN(Clk_r), .Q(Packet_Out[14]) );
  FDN1QM1P \Queue_reg[1][13]  ( .D(n426), .CPN(Clk_r), .Q(\Queue[1][13] ) );
  FDN1QM1P \Queue_reg[0][13]  ( .D(n458), .CPN(Clk_r), .Q(Packet_Out[13]) );
  FDN1QM1P \Queue_reg[1][12]  ( .D(n425), .CPN(Clk_r), .Q(\Queue[1][12] ) );
  FDN1QM1P \Queue_reg[0][12]  ( .D(n457), .CPN(Clk_r), .Q(Packet_Out[12]) );
  FDN1QM1P \Queue_reg[1][11]  ( .D(n424), .CPN(Clk_r), .Q(\Queue[1][11] ) );
  FDN1QM1P \Queue_reg[0][11]  ( .D(n456), .CPN(Clk_r), .Q(Packet_Out[11]) );
  FDN1QM1P \Queue_reg[1][10]  ( .D(n423), .CPN(Clk_r), .Q(\Queue[1][10] ) );
  FDN1QM1P \Queue_reg[0][10]  ( .D(n455), .CPN(Clk_r), .Q(Packet_Out[10]) );
  FDN1QM1P \Queue_reg[1][9]  ( .D(n422), .CPN(Clk_r), .Q(\Queue[1][9] ) );
  FDN1QM1P \Queue_reg[0][9]  ( .D(n454), .CPN(Clk_r), .Q(Packet_Out[9]) );
  FDN1QM1P \Queue_reg[1][8]  ( .D(n421), .CPN(Clk_r), .Q(\Queue[1][8] ) );
  FDN1QM1P \Queue_reg[0][8]  ( .D(n453), .CPN(Clk_r), .Q(Packet_Out[8]) );
  FDN1QM1P \Queue_reg[1][7]  ( .D(n420), .CPN(Clk_r), .Q(\Queue[1][7] ) );
  FDN1QM1P \Queue_reg[0][7]  ( .D(n452), .CPN(Clk_r), .Q(Packet_Out[7]) );
  FDN1QM1P \Queue_reg[1][6]  ( .D(n419), .CPN(Clk_r), .Q(\Queue[1][6] ) );
  FDN1QM1P \Queue_reg[0][6]  ( .D(n451), .CPN(Clk_r), .Q(Packet_Out[6]) );
  FDN1QM1P \Queue_reg[1][5]  ( .D(n418), .CPN(Clk_r), .Q(\Queue[1][5] ) );
  FDN1QM1P \Queue_reg[0][5]  ( .D(n450), .CPN(Clk_r), .Q(Packet_Out[5]) );
  FDN1QM1P \Queue_reg[1][4]  ( .D(n417), .CPN(Clk_r), .Q(\Queue[1][4] ) );
  FDN1QM1P \Queue_reg[0][4]  ( .D(n449), .CPN(Clk_r), .Q(Packet_Out[4]) );
  FDN1QM1P \Queue_reg[1][3]  ( .D(n416), .CPN(Clk_r), .Q(\Queue[1][3] ) );
  FDN1QM1P \Queue_reg[0][3]  ( .D(n448), .CPN(Clk_r), .Q(Packet_Out[3]) );
  FDN1QM1P \Queue_reg[1][2]  ( .D(n415), .CPN(Clk_r), .Q(\Queue[1][2] ) );
  FDN1QM1P \Queue_reg[0][2]  ( .D(n447), .CPN(Clk_r), .Q(Packet_Out[2]) );
  FDN1QM1P \Queue_reg[1][1]  ( .D(n414), .CPN(Clk_r), .Q(\Queue[1][1] ) );
  FDN1QM1P \Queue_reg[0][1]  ( .D(n446), .CPN(Clk_r), .Q(Packet_Out[1]) );
  FDN1QM1P \Queue_reg[1][0]  ( .D(n413), .CPN(Clk_r), .Q(\Queue[1][0] ) );
  FDN1QM1P \Queue_reg[0][0]  ( .D(n445), .CPN(Clk_r), .Q(Packet_Out[0]) );
  FDN2QM1P Empty_reg ( .D(n542), .CPN(Clk_r), .CD(Rst_n), .Q(n541) );
  BUFM2P U3 ( .A(n97), .Z(n7) );
  BUFM1P U4 ( .A(n97), .Z(n8) );
  BUFM1P U5 ( .A(n135), .Z(n10) );
  BUFM1P U6 ( .A(n135), .Z(n11) );
  BUFM1P U7 ( .A(n135), .Z(n12) );
  OAI211M4P U8 ( .A(n142), .B(n137), .C(Write_Ack), .D(n136), .Z(n208) );
  NR3M1P U9 ( .A(Count[2]), .B(n23), .C(n22), .Z(n140) );
  N1M1P U10 ( .A(Read_Ack), .Z(n137) );
  NR3M1P U11 ( .A(Count[0]), .B(Count[2]), .C(n22), .Z(n100) );
  N1M2P U12 ( .A(n18), .Z(n139) );
  OAI211M1P U13 ( .A(n140), .B(n137), .C(Write_Ack), .D(n98), .Z(n135) );
  NR3M1P U14 ( .A(n23), .B(Count[2]), .C(Count[1]), .Z(n376) );
  OAI211M4P U15 ( .A(n100), .B(n137), .C(Write_Ack), .D(n24), .Z(n59) );
  BUFM2P U16 ( .A(n132), .Z(n9) );
  BUFM2P U17 ( .A(n95), .Z(n6) );
  OAI21M2P U18 ( .A(Write_Ack), .B(Read_Ack), .C(n24), .Z(n56) );
  OAI211M4P U19 ( .A(n100), .B(n139), .C(Rst_n), .D(n138), .Z(n133) );
  NR2FM3P U20 ( .A(n61), .B(n21), .Z(n20) );
  OAI211M4P U21 ( .A(n140), .B(n139), .C(Rst_n), .D(n138), .Z(n206) );
  NR3M1P U22 ( .A(Count[0]), .B(Count[1]), .C(n19), .Z(n142) );
  AOI21M2P U23 ( .A(Write_Ack), .B(n100), .C(n141), .Z(n57) );
  N1M1P U24 ( .A(n142), .Z(n21) );
  N1M3P U25 ( .A(Write_Ack), .Z(n99) );
  N1M1P U26 ( .A(Count[0]), .Z(n23) );
  N1M1P U27 ( .A(Count[2]), .Z(n19) );
  N1M1P U28 ( .A(Count[1]), .Z(n22) );
  ND2M2P U29 ( .A(n18), .B(Rst_n), .Z(n61) );
  ND2M2P U30 ( .A(Read_Ack), .B(Rst_n), .Z(n141) );
  N1M1P U31 ( .A(Packet_In[2]), .Z(n148) );
  N1M1P U32 ( .A(Packet_In[6]), .Z(n156) );
  N1M1P U33 ( .A(Packet_In[7]), .Z(n158) );
  N1M1P U34 ( .A(Packet_In[3]), .Z(n150) );
  N1M1P U35 ( .A(Packet_In[5]), .Z(n154) );
  N1M1P U36 ( .A(Packet_In[4]), .Z(n152) );
  N1M1P U37 ( .A(Packet_In[8]), .Z(n160) );
  N1M1P U38 ( .A(Packet_In[0]), .Z(n144) );
  N1M1P U39 ( .A(Packet_In[10]), .Z(n164) );
  N1M1P U40 ( .A(Packet_In[11]), .Z(n166) );
  N1M1P U41 ( .A(Packet_In[9]), .Z(n162) );
  N1M1P U42 ( .A(Packet_In[20]), .Z(n184) );
  N1M1P U43 ( .A(Packet_In[14]), .Z(n172) );
  N1M1P U44 ( .A(Packet_In[13]), .Z(n170) );
  N1M1P U45 ( .A(Packet_In[27]), .Z(n198) );
  N1M1P U46 ( .A(Packet_In[23]), .Z(n190) );
  N1M1P U47 ( .A(Packet_In[25]), .Z(n194) );
  N1M1P U48 ( .A(Packet_In[1]), .Z(n146) );
  N1M1P U49 ( .A(Packet_In[29]), .Z(n202) );
  N1M1P U50 ( .A(Packet_In[22]), .Z(n188) );
  N1M1P U51 ( .A(Packet_In[28]), .Z(n200) );
  N1M1P U52 ( .A(Packet_In[19]), .Z(n182) );
  N1M1P U53 ( .A(Packet_In[21]), .Z(n186) );
  N1M1P U54 ( .A(Packet_In[18]), .Z(n180) );
  N1M1P U55 ( .A(Packet_In[12]), .Z(n168) );
  N1M1P U56 ( .A(Packet_In[26]), .Z(n196) );
  N1M1P U57 ( .A(Packet_In[17]), .Z(n178) );
  N1M1P U58 ( .A(Packet_In[16]), .Z(n176) );
  N1M1P U59 ( .A(Packet_In[24]), .Z(n192) );
  N1M1P U60 ( .A(Packet_In[15]), .Z(n174) );
  N1M1P U61 ( .A(Packet_In[31]), .Z(n373) );
  N1M1P U62 ( .A(Packet_In[30]), .Z(n204) );
  AOI21M6P U63 ( .A(Write_Ack), .B(n142), .C(n141), .Z(n205) );
  N1M2P U64 ( .A(n62), .Z(n94) );
  OAI211M1P U65 ( .A(n376), .B(n137), .C(Write_Ack), .D(n62), .Z(n97) );
  BUFM2P U66 ( .A(n56), .Z(n3) );
  BUFM2P U67 ( .A(n56), .Z(n4) );
  BUFM2P U68 ( .A(n57), .Z(n5) );
  NR2FM2P U69 ( .A(Read_Ack), .B(n99), .Z(n18) );
  AOI22M1P U70 ( .A(Count[0]), .B(n139), .C(n17), .D(n23), .Z(n14) );
  OA21M1P U71 ( .A(n139), .B(n100), .C(Rst_n), .Z(n98) );
  NR2M1P U72 ( .A(n137), .B(Write_Ack), .Z(n375) );
  NR2M1P U73 ( .A(n18), .B(n375), .Z(n374) );
  AOI22CDNM1P U74 ( .A(n374), .B(n23), .C(n374), .D(n23), .Z(n377) );
  N1M1P U75 ( .A(n375), .Z(n17) );
  AOI22CDNM1P U76 ( .A(Count[1]), .B(n14), .C(n14), .D(Count[1]), .Z(n378) );
  ND3M1P U77 ( .A(n23), .B(n19), .C(n22), .Z(n60) );
  ND2M1P U78 ( .A(Count[1]), .B(Read_Ack), .Z(n13) );
  OAI211M1P U79 ( .A(Count[1]), .B(n139), .C(n14), .D(n13), .Z(n15) );
  AOI22M1P U80 ( .A(n18), .B(n140), .C(Count[2]), .D(n15), .Z(n16) );
  OAI21M1P U81 ( .A(n60), .B(n17), .C(n16), .Z(n379) );
  AOI22CDNM1P U82 ( .A(n20), .B(n373), .C(\Queue[4][31] ), .D(n20), .Z(n380)
         );
  AOI22CDNM1P U83 ( .A(n20), .B(n144), .C(\Queue[4][0] ), .D(n20), .Z(n381) );
  AOI22CDNM1P U84 ( .A(n20), .B(n146), .C(\Queue[4][1] ), .D(n20), .Z(n382) );
  AOI22CDNM1P U85 ( .A(n20), .B(n148), .C(\Queue[4][2] ), .D(n20), .Z(n383) );
  AOI22CDNM1P U86 ( .A(n20), .B(n150), .C(\Queue[4][3] ), .D(n20), .Z(n384) );
  AOI22CDNM1P U87 ( .A(n20), .B(n152), .C(\Queue[4][4] ), .D(n20), .Z(n385) );
  AOI22CDNM1P U88 ( .A(n20), .B(n154), .C(\Queue[4][5] ), .D(n20), .Z(n386) );
  AOI22CDNM1P U89 ( .A(n20), .B(n156), .C(\Queue[4][6] ), .D(n20), .Z(n387) );
  AOI22CDNM1P U90 ( .A(n20), .B(n158), .C(\Queue[4][7] ), .D(n20), .Z(n388) );
  AOI22CDNM1P U91 ( .A(n20), .B(n160), .C(\Queue[4][8] ), .D(n20), .Z(n389) );
  AOI22CDNM1P U92 ( .A(n20), .B(n162), .C(\Queue[4][9] ), .D(n20), .Z(n390) );
  AOI22CDNM1P U93 ( .A(n20), .B(n164), .C(\Queue[4][10] ), .D(n20), .Z(n391)
         );
  AOI22CDNM1P U94 ( .A(n20), .B(n166), .C(\Queue[4][11] ), .D(n20), .Z(n392)
         );
  AOI22CDNM1P U95 ( .A(n20), .B(n168), .C(\Queue[4][12] ), .D(n20), .Z(n393)
         );
  AOI22CDNM1P U96 ( .A(n20), .B(n170), .C(\Queue[4][13] ), .D(n20), .Z(n394)
         );
  AOI22CDNM1P U97 ( .A(n20), .B(n172), .C(\Queue[4][14] ), .D(n20), .Z(n395)
         );
  AOI22CDNM1P U98 ( .A(n20), .B(n174), .C(\Queue[4][15] ), .D(n20), .Z(n396)
         );
  AOI22CDNM1P U99 ( .A(n20), .B(n176), .C(\Queue[4][16] ), .D(n20), .Z(n397)
         );
  AOI22CDNM1P U100 ( .A(n20), .B(n178), .C(\Queue[4][17] ), .D(n20), .Z(n398)
         );
  AOI22CDNM1P U101 ( .A(n20), .B(n180), .C(\Queue[4][18] ), .D(n20), .Z(n399)
         );
  AOI22CDNM1P U102 ( .A(n20), .B(n182), .C(\Queue[4][19] ), .D(n20), .Z(n400)
         );
  AOI22CDNM1P U103 ( .A(n20), .B(n184), .C(\Queue[4][20] ), .D(n20), .Z(n401)
         );
  AOI22CDNM1P U104 ( .A(n20), .B(n186), .C(\Queue[4][21] ), .D(n20), .Z(n402)
         );
  AOI22CDNM1P U105 ( .A(n20), .B(n188), .C(\Queue[4][22] ), .D(n20), .Z(n403)
         );
  AOI22CDNM1P U106 ( .A(n20), .B(n190), .C(\Queue[4][23] ), .D(n20), .Z(n404)
         );
  AOI22CDNM1P U107 ( .A(n20), .B(n192), .C(\Queue[4][24] ), .D(n20), .Z(n405)
         );
  AOI22CDNM1P U108 ( .A(n20), .B(n194), .C(\Queue[4][25] ), .D(n20), .Z(n406)
         );
  AOI22CDNM1P U109 ( .A(n20), .B(n196), .C(\Queue[4][26] ), .D(n20), .Z(n407)
         );
  AOI22CDNM1P U110 ( .A(n20), .B(n198), .C(\Queue[4][27] ), .D(n20), .Z(n408)
         );
  AOI22CDNM1P U111 ( .A(n20), .B(n200), .C(\Queue[4][28] ), .D(n20), .Z(n409)
         );
  AOI22CDNM1P U112 ( .A(n20), .B(n202), .C(\Queue[4][29] ), .D(n20), .Z(n410)
         );
  AOI22CDNM1P U113 ( .A(n20), .B(n204), .C(\Queue[4][30] ), .D(n20), .Z(n411)
         );
  OAI22CDNM1P U114 ( .A(n139), .B(n21), .C(n374), .D(Full), .Z(n412) );
  OA21M1P U115 ( .A(n139), .B(n376), .C(Rst_n), .Z(n24) );
  AOI22M1P U116 ( .A(\Queue[2][0] ), .B(n5), .C(\Queue[1][0] ), .D(n56), .Z(
        n25) );
  OAI21M1P U117 ( .A(n144), .B(n59), .C(n25), .Z(n413) );
  AOI22M1P U118 ( .A(n5), .B(\Queue[2][1] ), .C(\Queue[1][1] ), .D(n4), .Z(n26) );
  OAI21M1P U119 ( .A(n59), .B(n146), .C(n26), .Z(n414) );
  AOI22M1P U120 ( .A(n5), .B(\Queue[2][2] ), .C(\Queue[1][2] ), .D(n56), .Z(
        n27) );
  OAI21M1P U121 ( .A(n59), .B(n148), .C(n27), .Z(n415) );
  AOI22M1P U122 ( .A(n5), .B(\Queue[2][3] ), .C(\Queue[1][3] ), .D(n56), .Z(
        n28) );
  OAI21M1P U123 ( .A(n59), .B(n150), .C(n28), .Z(n416) );
  AOI22M1P U124 ( .A(n5), .B(\Queue[2][4] ), .C(\Queue[1][4] ), .D(n56), .Z(
        n29) );
  OAI21M1P U125 ( .A(n59), .B(n152), .C(n29), .Z(n417) );
  AOI22M1P U126 ( .A(n5), .B(\Queue[2][5] ), .C(\Queue[1][5] ), .D(n56), .Z(
        n30) );
  OAI21M1P U127 ( .A(n59), .B(n154), .C(n30), .Z(n418) );
  AOI22M1P U128 ( .A(n5), .B(\Queue[2][6] ), .C(\Queue[1][6] ), .D(n56), .Z(
        n31) );
  OAI21M1P U129 ( .A(n59), .B(n156), .C(n31), .Z(n419) );
  AOI22M1P U130 ( .A(n5), .B(\Queue[2][7] ), .C(\Queue[1][7] ), .D(n56), .Z(
        n32) );
  OAI21M1P U131 ( .A(n59), .B(n158), .C(n32), .Z(n420) );
  AOI22M1P U132 ( .A(n5), .B(\Queue[2][8] ), .C(\Queue[1][8] ), .D(n56), .Z(
        n33) );
  OAI21M1P U133 ( .A(n59), .B(n160), .C(n33), .Z(n421) );
  AOI22M1P U134 ( .A(n5), .B(\Queue[2][9] ), .C(\Queue[1][9] ), .D(n3), .Z(n34) );
  OAI21M1P U135 ( .A(n59), .B(n162), .C(n34), .Z(n422) );
  AOI22M1P U136 ( .A(n5), .B(\Queue[2][10] ), .C(\Queue[1][10] ), .D(n3), .Z(
        n35) );
  OAI21M1P U137 ( .A(n59), .B(n164), .C(n35), .Z(n423) );
  AOI22M1P U138 ( .A(n5), .B(\Queue[2][11] ), .C(\Queue[1][11] ), .D(n3), .Z(
        n36) );
  OAI21M1P U139 ( .A(n59), .B(n166), .C(n36), .Z(n424) );
  AOI22M1P U140 ( .A(n57), .B(\Queue[2][12] ), .C(\Queue[1][12] ), .D(n3), .Z(
        n37) );
  OAI21M1P U141 ( .A(n59), .B(n168), .C(n37), .Z(n425) );
  AOI22M1P U142 ( .A(n57), .B(\Queue[2][13] ), .C(\Queue[1][13] ), .D(n3), .Z(
        n38) );
  OAI21M1P U143 ( .A(n59), .B(n170), .C(n38), .Z(n426) );
  AOI22M1P U144 ( .A(n57), .B(\Queue[2][14] ), .C(\Queue[1][14] ), .D(n3), .Z(
        n39) );
  OAI21M1P U145 ( .A(n59), .B(n172), .C(n39), .Z(n427) );
  AOI22M1P U146 ( .A(n57), .B(\Queue[2][15] ), .C(\Queue[1][15] ), .D(n3), .Z(
        n40) );
  OAI21M1P U147 ( .A(n59), .B(n174), .C(n40), .Z(n428) );
  AOI22M1P U148 ( .A(n57), .B(\Queue[2][16] ), .C(\Queue[1][16] ), .D(n3), .Z(
        n41) );
  OAI21M1P U149 ( .A(n59), .B(n176), .C(n41), .Z(n429) );
  AOI22M1P U150 ( .A(n57), .B(\Queue[2][17] ), .C(\Queue[1][17] ), .D(n3), .Z(
        n42) );
  OAI21M1P U151 ( .A(n59), .B(n178), .C(n42), .Z(n430) );
  AOI22M1P U152 ( .A(n57), .B(\Queue[2][18] ), .C(\Queue[1][18] ), .D(n4), .Z(
        n43) );
  OAI21M1P U153 ( .A(n59), .B(n180), .C(n43), .Z(n431) );
  AOI22M1P U154 ( .A(n57), .B(\Queue[2][19] ), .C(\Queue[1][19] ), .D(n4), .Z(
        n44) );
  OAI21M1P U155 ( .A(n59), .B(n182), .C(n44), .Z(n432) );
  AOI22M1P U156 ( .A(n57), .B(\Queue[2][20] ), .C(\Queue[1][20] ), .D(n4), .Z(
        n45) );
  OAI21M1P U157 ( .A(n59), .B(n184), .C(n45), .Z(n433) );
  AOI22M1P U158 ( .A(n57), .B(\Queue[2][21] ), .C(\Queue[1][21] ), .D(n4), .Z(
        n46) );
  OAI21M1P U159 ( .A(n59), .B(n186), .C(n46), .Z(n434) );
  AOI22M1P U160 ( .A(n5), .B(\Queue[2][22] ), .C(\Queue[1][22] ), .D(n4), .Z(
        n47) );
  OAI21M1P U161 ( .A(n59), .B(n188), .C(n47), .Z(n435) );
  AOI22M1P U162 ( .A(n5), .B(\Queue[2][23] ), .C(\Queue[1][23] ), .D(n4), .Z(
        n48) );
  OAI21M1P U163 ( .A(n59), .B(n190), .C(n48), .Z(n436) );
  AOI22M1P U164 ( .A(n5), .B(\Queue[2][24] ), .C(\Queue[1][24] ), .D(n4), .Z(
        n49) );
  OAI21M1P U165 ( .A(n59), .B(n192), .C(n49), .Z(n437) );
  AOI22M1P U166 ( .A(n57), .B(\Queue[2][25] ), .C(\Queue[1][25] ), .D(n4), .Z(
        n50) );
  OAI21M1P U167 ( .A(n59), .B(n194), .C(n50), .Z(n438) );
  AOI22M1P U168 ( .A(n57), .B(\Queue[2][26] ), .C(\Queue[1][26] ), .D(n4), .Z(
        n51) );
  OAI21M1P U169 ( .A(n59), .B(n196), .C(n51), .Z(n439) );
  AOI22M1P U170 ( .A(n57), .B(\Queue[2][27] ), .C(\Queue[1][27] ), .D(n3), .Z(
        n52) );
  OAI21M1P U171 ( .A(n59), .B(n198), .C(n52), .Z(n440) );
  AOI22M1P U172 ( .A(n57), .B(\Queue[2][28] ), .C(\Queue[1][28] ), .D(n4), .Z(
        n53) );
  OAI21M1P U173 ( .A(n59), .B(n200), .C(n53), .Z(n441) );
  AOI22M1P U174 ( .A(n57), .B(\Queue[2][29] ), .C(\Queue[1][29] ), .D(n3), .Z(
        n54) );
  OAI21M1P U175 ( .A(n59), .B(n202), .C(n54), .Z(n442) );
  AOI22M1P U176 ( .A(n57), .B(\Queue[2][30] ), .C(\Queue[1][30] ), .D(n3), .Z(
        n55) );
  OAI21M1P U177 ( .A(n59), .B(n204), .C(n55), .Z(n443) );
  AOI22M1P U178 ( .A(n57), .B(\Queue[2][31] ), .C(\Queue[1][31] ), .D(n4), .Z(
        n58) );
  OAI21M1P U179 ( .A(n59), .B(n373), .C(n58), .Z(n444) );
  OAI21M1P U180 ( .A(n61), .B(n60), .C(n141), .Z(n62) );
  AOI21M1P U181 ( .A(Write_Ack), .B(n376), .C(n141), .Z(n95) );
  AOI22M1P U182 ( .A(\Queue[1][0] ), .B(n6), .C(n94), .D(Packet_Out[0]), .Z(
        n63) );
  OAI21M1P U183 ( .A(n144), .B(n7), .C(n63), .Z(n445) );
  AOI22M1P U184 ( .A(\Queue[1][1] ), .B(n6), .C(n94), .D(Packet_Out[1]), .Z(
        n64) );
  OAI21M1P U185 ( .A(n146), .B(n7), .C(n64), .Z(n446) );
  AOI22M1P U186 ( .A(\Queue[1][2] ), .B(n6), .C(n94), .D(Packet_Out[2]), .Z(
        n65) );
  OAI21M1P U187 ( .A(n148), .B(n7), .C(n65), .Z(n447) );
  AOI22M1P U188 ( .A(\Queue[1][3] ), .B(n6), .C(n94), .D(Packet_Out[3]), .Z(
        n66) );
  OAI21M1P U189 ( .A(n150), .B(n7), .C(n66), .Z(n448) );
  AOI22M1P U190 ( .A(\Queue[1][4] ), .B(n6), .C(n94), .D(Packet_Out[4]), .Z(
        n67) );
  OAI21M1P U191 ( .A(n152), .B(n7), .C(n67), .Z(n449) );
  AOI22M1P U192 ( .A(\Queue[1][5] ), .B(n6), .C(n94), .D(Packet_Out[5]), .Z(
        n68) );
  OAI21M1P U193 ( .A(n154), .B(n7), .C(n68), .Z(n450) );
  AOI22M1P U194 ( .A(\Queue[1][6] ), .B(n6), .C(n94), .D(Packet_Out[6]), .Z(
        n69) );
  OAI21M1P U195 ( .A(n156), .B(n7), .C(n69), .Z(n451) );
  AOI22M1P U196 ( .A(\Queue[1][7] ), .B(n6), .C(n94), .D(Packet_Out[7]), .Z(
        n70) );
  OAI21M1P U197 ( .A(n158), .B(n7), .C(n70), .Z(n452) );
  AOI22M1P U198 ( .A(\Queue[1][8] ), .B(n6), .C(n94), .D(Packet_Out[8]), .Z(
        n71) );
  OAI21M1P U199 ( .A(n160), .B(n7), .C(n71), .Z(n453) );
  AOI22M1P U200 ( .A(\Queue[1][9] ), .B(n6), .C(n94), .D(Packet_Out[9]), .Z(
        n72) );
  OAI21M1P U201 ( .A(n162), .B(n7), .C(n72), .Z(n454) );
  AOI22M1P U202 ( .A(\Queue[1][10] ), .B(n95), .C(n94), .D(Packet_Out[10]), 
        .Z(n73) );
  OAI21M1P U203 ( .A(n164), .B(n7), .C(n73), .Z(n455) );
  AOI22M1P U204 ( .A(\Queue[1][11] ), .B(n95), .C(n94), .D(Packet_Out[11]), 
        .Z(n74) );
  OAI21M1P U205 ( .A(n166), .B(n7), .C(n74), .Z(n456) );
  AOI22M1P U206 ( .A(\Queue[1][12] ), .B(n95), .C(n94), .D(Packet_Out[12]), 
        .Z(n75) );
  OAI21M1P U207 ( .A(n168), .B(n7), .C(n75), .Z(n457) );
  AOI22M1P U208 ( .A(\Queue[1][13] ), .B(n95), .C(n94), .D(Packet_Out[13]), 
        .Z(n76) );
  OAI21M1P U209 ( .A(n170), .B(n7), .C(n76), .Z(n458) );
  AOI22M1P U210 ( .A(\Queue[1][14] ), .B(n95), .C(n94), .D(Packet_Out[14]), 
        .Z(n77) );
  OAI21M1P U211 ( .A(n172), .B(n7), .C(n77), .Z(n459) );
  AOI22M1P U212 ( .A(\Queue[1][15] ), .B(n95), .C(n94), .D(Packet_Out[15]), 
        .Z(n78) );
  OAI21M1P U213 ( .A(n174), .B(n7), .C(n78), .Z(n460) );
  AOI22M1P U214 ( .A(\Queue[1][16] ), .B(n6), .C(n94), .D(Packet_Out[16]), .Z(
        n79) );
  OAI21M1P U215 ( .A(n176), .B(n7), .C(n79), .Z(n461) );
  AOI22M1P U216 ( .A(\Queue[1][17] ), .B(n6), .C(n94), .D(Packet_Out[17]), .Z(
        n80) );
  OAI21M1P U217 ( .A(n178), .B(n7), .C(n80), .Z(n462) );
  AOI22M1P U218 ( .A(\Queue[1][18] ), .B(n6), .C(n94), .D(Packet_Out[18]), .Z(
        n81) );
  OAI21M1P U219 ( .A(n180), .B(n7), .C(n81), .Z(n463) );
  AOI22M1P U220 ( .A(\Queue[1][19] ), .B(n6), .C(n94), .D(Packet_Out[19]), .Z(
        n82) );
  OAI21M1P U221 ( .A(n182), .B(n7), .C(n82), .Z(n464) );
  AOI22M1P U222 ( .A(\Queue[1][20] ), .B(n6), .C(n94), .D(Packet_Out[20]), .Z(
        n83) );
  OAI21M1P U223 ( .A(n184), .B(n8), .C(n83), .Z(n465) );
  AOI22M1P U224 ( .A(\Queue[1][21] ), .B(n6), .C(n94), .D(Packet_Out[21]), .Z(
        n84) );
  OAI21M1P U225 ( .A(n186), .B(n8), .C(n84), .Z(n466) );
  AOI22M1P U226 ( .A(\Queue[1][22] ), .B(n6), .C(n94), .D(Packet_Out[22]), .Z(
        n85) );
  OAI21M1P U227 ( .A(n188), .B(n8), .C(n85), .Z(n467) );
  AOI22M1P U228 ( .A(\Queue[1][23] ), .B(n6), .C(n94), .D(Packet_Out[23]), .Z(
        n86) );
  OAI21M1P U229 ( .A(n190), .B(n8), .C(n86), .Z(n468) );
  AOI22M1P U230 ( .A(\Queue[1][24] ), .B(n6), .C(n94), .D(Packet_Out[24]), .Z(
        n87) );
  OAI21M1P U231 ( .A(n192), .B(n8), .C(n87), .Z(n469) );
  AOI22M1P U232 ( .A(\Queue[1][25] ), .B(n6), .C(n94), .D(Packet_Out[25]), .Z(
        n88) );
  OAI21M1P U233 ( .A(n194), .B(n8), .C(n88), .Z(n470) );
  AOI22M1P U234 ( .A(\Queue[1][26] ), .B(n6), .C(n94), .D(Packet_Out[26]), .Z(
        n89) );
  OAI21M1P U235 ( .A(n196), .B(n8), .C(n89), .Z(n471) );
  AOI22M1P U236 ( .A(\Queue[1][27] ), .B(n6), .C(n94), .D(Packet_Out[27]), .Z(
        n90) );
  OAI21M1P U237 ( .A(n198), .B(n8), .C(n90), .Z(n472) );
  AOI22M1P U238 ( .A(\Queue[1][28] ), .B(n6), .C(n94), .D(Packet_Out[28]), .Z(
        n91) );
  OAI21M1P U239 ( .A(n200), .B(n8), .C(n91), .Z(n473) );
  AOI22M1P U240 ( .A(\Queue[1][29] ), .B(n6), .C(n94), .D(Packet_Out[29]), .Z(
        n92) );
  OAI21M1P U241 ( .A(n202), .B(n8), .C(n92), .Z(n474) );
  AOI22M1P U242 ( .A(\Queue[1][30] ), .B(n6), .C(n94), .D(Packet_Out[30]), .Z(
        n93) );
  OAI21M1P U243 ( .A(n204), .B(n7), .C(n93), .Z(n475) );
  AOI22M1P U244 ( .A(\Queue[1][31] ), .B(n6), .C(n94), .D(Packet_Out[31]), .Z(
        n96) );
  OAI21M1P U245 ( .A(n373), .B(n8), .C(n96), .Z(n476) );
  ND2M1P U246 ( .A(n99), .B(n137), .Z(n138) );
  AOI21M1P U247 ( .A(Write_Ack), .B(n140), .C(n141), .Z(n132) );
  AOI22M1P U248 ( .A(\Queue[2][0] ), .B(n133), .C(\Queue[3][0] ), .D(n132), 
        .Z(n101) );
  OAI21M1P U249 ( .A(n144), .B(n10), .C(n101), .Z(n477) );
  AOI22M1P U250 ( .A(\Queue[2][1] ), .B(n133), .C(n9), .D(\Queue[3][1] ), .Z(
        n102) );
  OAI21M1P U251 ( .A(n146), .B(n10), .C(n102), .Z(n478) );
  AOI22M1P U252 ( .A(\Queue[2][2] ), .B(n133), .C(n9), .D(\Queue[3][2] ), .Z(
        n103) );
  OAI21M1P U253 ( .A(n148), .B(n10), .C(n103), .Z(n479) );
  AOI22M1P U254 ( .A(\Queue[2][3] ), .B(n133), .C(n9), .D(\Queue[3][3] ), .Z(
        n104) );
  OAI21M1P U255 ( .A(n150), .B(n10), .C(n104), .Z(n480) );
  AOI22M1P U256 ( .A(\Queue[2][4] ), .B(n133), .C(n9), .D(\Queue[3][4] ), .Z(
        n105) );
  OAI21M1P U257 ( .A(n152), .B(n10), .C(n105), .Z(n481) );
  AOI22M1P U258 ( .A(\Queue[2][5] ), .B(n133), .C(n9), .D(\Queue[3][5] ), .Z(
        n106) );
  OAI21M1P U259 ( .A(n154), .B(n10), .C(n106), .Z(n482) );
  AOI22M1P U260 ( .A(\Queue[2][6] ), .B(n133), .C(n9), .D(\Queue[3][6] ), .Z(
        n107) );
  OAI21M1P U261 ( .A(n156), .B(n10), .C(n107), .Z(n483) );
  AOI22M1P U262 ( .A(\Queue[2][7] ), .B(n133), .C(n132), .D(\Queue[3][7] ), 
        .Z(n108) );
  OAI21M1P U263 ( .A(n158), .B(n10), .C(n108), .Z(n484) );
  AOI22M1P U264 ( .A(\Queue[2][8] ), .B(n133), .C(n132), .D(\Queue[3][8] ), 
        .Z(n109) );
  OAI21M1P U265 ( .A(n160), .B(n10), .C(n109), .Z(n485) );
  AOI22M1P U266 ( .A(\Queue[2][9] ), .B(n133), .C(n132), .D(\Queue[3][9] ), 
        .Z(n110) );
  OAI21M1P U267 ( .A(n162), .B(n10), .C(n110), .Z(n486) );
  AOI22M1P U268 ( .A(\Queue[2][10] ), .B(n133), .C(n132), .D(\Queue[3][10] ), 
        .Z(n111) );
  OAI21M1P U269 ( .A(n164), .B(n11), .C(n111), .Z(n487) );
  AOI22M1P U270 ( .A(\Queue[2][11] ), .B(n133), .C(n132), .D(\Queue[3][11] ), 
        .Z(n112) );
  OAI21M1P U271 ( .A(n166), .B(n11), .C(n112), .Z(n488) );
  AOI22M1P U272 ( .A(\Queue[2][12] ), .B(n133), .C(n9), .D(\Queue[3][12] ), 
        .Z(n113) );
  OAI21M1P U273 ( .A(n168), .B(n11), .C(n113), .Z(n489) );
  AOI22M1P U274 ( .A(\Queue[2][13] ), .B(n133), .C(n9), .D(\Queue[3][13] ), 
        .Z(n114) );
  OAI21M1P U275 ( .A(n170), .B(n11), .C(n114), .Z(n490) );
  AOI22M1P U276 ( .A(\Queue[2][14] ), .B(n133), .C(n9), .D(\Queue[3][14] ), 
        .Z(n115) );
  OAI21M1P U277 ( .A(n172), .B(n11), .C(n115), .Z(n491) );
  AOI22M1P U278 ( .A(\Queue[2][15] ), .B(n133), .C(n9), .D(\Queue[3][15] ), 
        .Z(n116) );
  OAI21M1P U279 ( .A(n174), .B(n11), .C(n116), .Z(n492) );
  AOI22M1P U280 ( .A(\Queue[2][16] ), .B(n133), .C(n9), .D(\Queue[3][16] ), 
        .Z(n117) );
  OAI21M1P U281 ( .A(n176), .B(n11), .C(n117), .Z(n493) );
  AOI22M1P U282 ( .A(\Queue[2][17] ), .B(n133), .C(n9), .D(\Queue[3][17] ), 
        .Z(n118) );
  OAI21M1P U283 ( .A(n178), .B(n11), .C(n118), .Z(n494) );
  AOI22M1P U284 ( .A(\Queue[2][18] ), .B(n133), .C(n9), .D(\Queue[3][18] ), 
        .Z(n119) );
  OAI21M1P U285 ( .A(n180), .B(n11), .C(n119), .Z(n495) );
  AOI22M1P U286 ( .A(\Queue[2][19] ), .B(n133), .C(n9), .D(\Queue[3][19] ), 
        .Z(n120) );
  OAI21M1P U287 ( .A(n182), .B(n11), .C(n120), .Z(n496) );
  AOI22M1P U288 ( .A(\Queue[2][20] ), .B(n133), .C(n9), .D(\Queue[3][20] ), 
        .Z(n121) );
  OAI21M1P U289 ( .A(n184), .B(n12), .C(n121), .Z(n497) );
  AOI22M1P U290 ( .A(\Queue[2][21] ), .B(n133), .C(n9), .D(\Queue[3][21] ), 
        .Z(n122) );
  OAI21M1P U291 ( .A(n186), .B(n12), .C(n122), .Z(n498) );
  AOI22M1P U292 ( .A(\Queue[2][22] ), .B(n133), .C(n9), .D(\Queue[3][22] ), 
        .Z(n123) );
  OAI21M1P U293 ( .A(n188), .B(n12), .C(n123), .Z(n499) );
  AOI22M1P U294 ( .A(\Queue[2][23] ), .B(n133), .C(n9), .D(\Queue[3][23] ), 
        .Z(n124) );
  OAI21M1P U295 ( .A(n190), .B(n12), .C(n124), .Z(n500) );
  AOI22M1P U296 ( .A(\Queue[2][24] ), .B(n133), .C(n9), .D(\Queue[3][24] ), 
        .Z(n125) );
  OAI21M1P U297 ( .A(n192), .B(n12), .C(n125), .Z(n501) );
  AOI22M1P U298 ( .A(\Queue[2][25] ), .B(n133), .C(n9), .D(\Queue[3][25] ), 
        .Z(n126) );
  OAI21M1P U299 ( .A(n194), .B(n12), .C(n126), .Z(n502) );
  AOI22M1P U300 ( .A(\Queue[2][26] ), .B(n133), .C(n9), .D(\Queue[3][26] ), 
        .Z(n127) );
  OAI21M1P U301 ( .A(n196), .B(n12), .C(n127), .Z(n503) );
  AOI22M1P U302 ( .A(\Queue[2][27] ), .B(n133), .C(n9), .D(\Queue[3][27] ), 
        .Z(n128) );
  OAI21M1P U303 ( .A(n198), .B(n12), .C(n128), .Z(n504) );
  AOI22M1P U304 ( .A(\Queue[2][28] ), .B(n133), .C(n9), .D(\Queue[3][28] ), 
        .Z(n129) );
  OAI21M1P U305 ( .A(n200), .B(n12), .C(n129), .Z(n505) );
  AOI22M1P U306 ( .A(\Queue[2][29] ), .B(n133), .C(n9), .D(\Queue[3][29] ), 
        .Z(n130) );
  OAI21M1P U307 ( .A(n202), .B(n12), .C(n130), .Z(n506) );
  AOI22M1P U308 ( .A(\Queue[2][30] ), .B(n133), .C(n9), .D(\Queue[3][30] ), 
        .Z(n131) );
  OAI21M1P U309 ( .A(n204), .B(n135), .C(n131), .Z(n507) );
  AOI22M1P U310 ( .A(\Queue[2][31] ), .B(n133), .C(n9), .D(\Queue[3][31] ), 
        .Z(n134) );
  OAI21M1P U311 ( .A(n373), .B(n135), .C(n134), .Z(n508) );
  OA21M1P U312 ( .A(n139), .B(n140), .C(Rst_n), .Z(n136) );
  AOI22M1P U313 ( .A(\Queue[3][0] ), .B(n206), .C(n205), .D(\Queue[4][0] ), 
        .Z(n143) );
  OAI21M1P U314 ( .A(n144), .B(n208), .C(n143), .Z(n509) );
  AOI22M1P U315 ( .A(\Queue[3][1] ), .B(n206), .C(n205), .D(\Queue[4][1] ), 
        .Z(n145) );
  OAI21M1P U316 ( .A(n146), .B(n208), .C(n145), .Z(n510) );
  AOI22M1P U317 ( .A(\Queue[3][2] ), .B(n206), .C(n205), .D(\Queue[4][2] ), 
        .Z(n147) );
  OAI21M1P U318 ( .A(n148), .B(n208), .C(n147), .Z(n511) );
  AOI22M1P U319 ( .A(\Queue[3][3] ), .B(n206), .C(n205), .D(\Queue[4][3] ), 
        .Z(n149) );
  OAI21M1P U320 ( .A(n150), .B(n208), .C(n149), .Z(n512) );
  AOI22M1P U321 ( .A(\Queue[3][4] ), .B(n206), .C(n205), .D(\Queue[4][4] ), 
        .Z(n151) );
  OAI21M1P U322 ( .A(n152), .B(n208), .C(n151), .Z(n513) );
  AOI22M1P U323 ( .A(\Queue[3][5] ), .B(n206), .C(n205), .D(\Queue[4][5] ), 
        .Z(n153) );
  OAI21M1P U324 ( .A(n154), .B(n208), .C(n153), .Z(n514) );
  AOI22M1P U325 ( .A(\Queue[3][6] ), .B(n206), .C(n205), .D(\Queue[4][6] ), 
        .Z(n155) );
  OAI21M1P U326 ( .A(n156), .B(n208), .C(n155), .Z(n515) );
  AOI22M1P U327 ( .A(\Queue[3][7] ), .B(n206), .C(n205), .D(\Queue[4][7] ), 
        .Z(n157) );
  OAI21M1P U328 ( .A(n158), .B(n208), .C(n157), .Z(n516) );
  AOI22M1P U329 ( .A(\Queue[3][8] ), .B(n206), .C(n205), .D(\Queue[4][8] ), 
        .Z(n159) );
  OAI21M1P U330 ( .A(n160), .B(n208), .C(n159), .Z(n517) );
  AOI22M1P U331 ( .A(\Queue[3][9] ), .B(n206), .C(n205), .D(\Queue[4][9] ), 
        .Z(n161) );
  OAI21M1P U332 ( .A(n162), .B(n208), .C(n161), .Z(n518) );
  AOI22M1P U333 ( .A(\Queue[3][10] ), .B(n206), .C(n205), .D(\Queue[4][10] ), 
        .Z(n163) );
  OAI21M1P U334 ( .A(n164), .B(n208), .C(n163), .Z(n519) );
  AOI22M1P U335 ( .A(\Queue[3][11] ), .B(n206), .C(n205), .D(\Queue[4][11] ), 
        .Z(n165) );
  OAI21M1P U336 ( .A(n166), .B(n208), .C(n165), .Z(n520) );
  AOI22M1P U337 ( .A(\Queue[3][12] ), .B(n206), .C(n205), .D(\Queue[4][12] ), 
        .Z(n167) );
  OAI21M1P U338 ( .A(n168), .B(n208), .C(n167), .Z(n521) );
  AOI22M1P U339 ( .A(\Queue[3][13] ), .B(n206), .C(n205), .D(\Queue[4][13] ), 
        .Z(n169) );
  OAI21M1P U340 ( .A(n170), .B(n208), .C(n169), .Z(n522) );
  AOI22M1P U341 ( .A(\Queue[3][14] ), .B(n206), .C(n205), .D(\Queue[4][14] ), 
        .Z(n171) );
  OAI21M1P U342 ( .A(n172), .B(n208), .C(n171), .Z(n523) );
  AOI22M1P U343 ( .A(\Queue[3][15] ), .B(n206), .C(n205), .D(\Queue[4][15] ), 
        .Z(n173) );
  OAI21M1P U344 ( .A(n174), .B(n208), .C(n173), .Z(n524) );
  AOI22M1P U345 ( .A(\Queue[3][16] ), .B(n206), .C(n205), .D(\Queue[4][16] ), 
        .Z(n175) );
  OAI21M1P U346 ( .A(n176), .B(n208), .C(n175), .Z(n525) );
  AOI22M1P U347 ( .A(\Queue[3][17] ), .B(n206), .C(n205), .D(\Queue[4][17] ), 
        .Z(n177) );
  OAI21M1P U348 ( .A(n178), .B(n208), .C(n177), .Z(n526) );
  AOI22M1P U349 ( .A(\Queue[3][18] ), .B(n206), .C(n205), .D(\Queue[4][18] ), 
        .Z(n179) );
  OAI21M1P U350 ( .A(n180), .B(n208), .C(n179), .Z(n527) );
  AOI22M1P U351 ( .A(\Queue[3][19] ), .B(n206), .C(n205), .D(\Queue[4][19] ), 
        .Z(n181) );
  OAI21M1P U352 ( .A(n182), .B(n208), .C(n181), .Z(n528) );
  AOI22M1P U353 ( .A(\Queue[3][20] ), .B(n206), .C(n205), .D(\Queue[4][20] ), 
        .Z(n183) );
  OAI21M1P U354 ( .A(n184), .B(n208), .C(n183), .Z(n529) );
  AOI22M1P U355 ( .A(\Queue[3][21] ), .B(n206), .C(n205), .D(\Queue[4][21] ), 
        .Z(n185) );
  OAI21M1P U356 ( .A(n186), .B(n208), .C(n185), .Z(n530) );
  AOI22M1P U357 ( .A(\Queue[3][22] ), .B(n206), .C(n205), .D(\Queue[4][22] ), 
        .Z(n187) );
  OAI21M1P U358 ( .A(n188), .B(n208), .C(n187), .Z(n531) );
  AOI22M1P U359 ( .A(\Queue[3][23] ), .B(n206), .C(n205), .D(\Queue[4][23] ), 
        .Z(n189) );
  OAI21M1P U360 ( .A(n190), .B(n208), .C(n189), .Z(n532) );
  AOI22M1P U361 ( .A(\Queue[3][24] ), .B(n206), .C(n205), .D(\Queue[4][24] ), 
        .Z(n191) );
  OAI21M1P U362 ( .A(n192), .B(n208), .C(n191), .Z(n533) );
  AOI22M1P U363 ( .A(\Queue[3][25] ), .B(n206), .C(n205), .D(\Queue[4][25] ), 
        .Z(n193) );
  OAI21M1P U364 ( .A(n194), .B(n208), .C(n193), .Z(n534) );
  AOI22M1P U365 ( .A(\Queue[3][26] ), .B(n206), .C(n205), .D(\Queue[4][26] ), 
        .Z(n195) );
  OAI21M1P U366 ( .A(n196), .B(n208), .C(n195), .Z(n535) );
  AOI22M1P U367 ( .A(\Queue[3][27] ), .B(n206), .C(n205), .D(\Queue[4][27] ), 
        .Z(n197) );
  OAI21M1P U368 ( .A(n198), .B(n208), .C(n197), .Z(n536) );
  AOI22M1P U369 ( .A(\Queue[3][28] ), .B(n206), .C(n205), .D(\Queue[4][28] ), 
        .Z(n199) );
  OAI21M1P U370 ( .A(n200), .B(n208), .C(n199), .Z(n537) );
  AOI22M1P U371 ( .A(\Queue[3][29] ), .B(n206), .C(n205), .D(\Queue[4][29] ), 
        .Z(n201) );
  OAI21M1P U372 ( .A(n202), .B(n208), .C(n201), .Z(n538) );
  AOI22M1P U373 ( .A(\Queue[3][30] ), .B(n206), .C(n205), .D(\Queue[4][30] ), 
        .Z(n203) );
  OAI21M1P U374 ( .A(n204), .B(n208), .C(n203), .Z(n539) );
  AOI22M1P U375 ( .A(\Queue[3][31] ), .B(n206), .C(n205), .D(\Queue[4][31] ), 
        .Z(n207) );
  OAI21M1P U376 ( .A(n373), .B(n208), .C(n207), .Z(n540) );
  N1M1P U377 ( .A(n541), .Z(Empty) );
  AOI22M1P U378 ( .A(n376), .B(n375), .C(n374), .D(Empty), .Z(n542) );
endmodule


module Packet_Queue_4 ( Clk_r, Rst_n, Packet_In, Read_Ack, Write_Ack, 
        Packet_Out, Empty, Full );
  input [31:0] Packet_In;
  output [31:0] Packet_Out;
  input Clk_r, Rst_n, Read_Ack, Write_Ack;
  output Empty, Full;
  wire   \Queue[4][31] , \Queue[4][30] , \Queue[4][29] , \Queue[4][28] ,
         \Queue[4][27] , \Queue[4][26] , \Queue[4][25] , \Queue[4][24] ,
         \Queue[4][23] , \Queue[4][22] , \Queue[4][21] , \Queue[4][20] ,
         \Queue[4][19] , \Queue[4][18] , \Queue[4][17] , \Queue[4][16] ,
         \Queue[4][15] , \Queue[4][14] , \Queue[4][13] , \Queue[4][12] ,
         \Queue[4][11] , \Queue[4][10] , \Queue[4][9] , \Queue[4][8] ,
         \Queue[4][7] , \Queue[4][6] , \Queue[4][5] , \Queue[4][4] ,
         \Queue[4][3] , \Queue[4][2] , \Queue[4][1] , \Queue[4][0] ,
         \Queue[3][31] , \Queue[3][30] , \Queue[3][29] , \Queue[3][28] ,
         \Queue[3][27] , \Queue[3][26] , \Queue[3][25] , \Queue[3][24] ,
         \Queue[3][23] , \Queue[3][22] , \Queue[3][21] , \Queue[3][20] ,
         \Queue[3][19] , \Queue[3][18] , \Queue[3][17] , \Queue[3][16] ,
         \Queue[3][15] , \Queue[3][14] , \Queue[3][13] , \Queue[3][12] ,
         \Queue[3][11] , \Queue[3][10] , \Queue[3][9] , \Queue[3][8] ,
         \Queue[3][7] , \Queue[3][6] , \Queue[3][5] , \Queue[3][4] ,
         \Queue[3][3] , \Queue[3][2] , \Queue[3][1] , \Queue[3][0] ,
         \Queue[2][31] , \Queue[2][30] , \Queue[2][29] , \Queue[2][28] ,
         \Queue[2][27] , \Queue[2][26] , \Queue[2][25] , \Queue[2][24] ,
         \Queue[2][23] , \Queue[2][22] , \Queue[2][21] , \Queue[2][20] ,
         \Queue[2][19] , \Queue[2][18] , \Queue[2][17] , \Queue[2][16] ,
         \Queue[2][15] , \Queue[2][14] , \Queue[2][13] , \Queue[2][12] ,
         \Queue[2][11] , \Queue[2][10] , \Queue[2][9] , \Queue[2][8] ,
         \Queue[2][7] , \Queue[2][6] , \Queue[2][5] , \Queue[2][4] ,
         \Queue[2][3] , \Queue[2][2] , \Queue[2][1] , \Queue[2][0] ,
         \Queue[1][31] , \Queue[1][30] , \Queue[1][29] , \Queue[1][28] ,
         \Queue[1][27] , \Queue[1][26] , \Queue[1][25] , \Queue[1][24] ,
         \Queue[1][23] , \Queue[1][22] , \Queue[1][21] , \Queue[1][20] ,
         \Queue[1][19] , \Queue[1][18] , \Queue[1][17] , \Queue[1][16] ,
         \Queue[1][15] , \Queue[1][14] , \Queue[1][13] , \Queue[1][12] ,
         \Queue[1][11] , \Queue[1][10] , \Queue[1][9] , \Queue[1][8] ,
         \Queue[1][7] , \Queue[1][6] , \Queue[1][5] , \Queue[1][4] ,
         \Queue[1][3] , \Queue[1][2] , \Queue[1][1] , \Queue[1][0] , n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541;
  wire   [2:0] Count;

  FDN2QM1P \Count_reg[0]  ( .D(n376), .CPN(Clk_r), .CD(Rst_n), .Q(Count[0]) );
  FDN2QM1P \Count_reg[1]  ( .D(n377), .CPN(Clk_r), .CD(Rst_n), .Q(Count[1]) );
  FDN2QM1P \Count_reg[2]  ( .D(n378), .CPN(Clk_r), .CD(Rst_n), .Q(Count[2]) );
  FDN1QM1P \Queue_reg[4][30]  ( .D(n410), .CPN(Clk_r), .Q(\Queue[4][30] ) );
  FDN1QM1P \Queue_reg[3][30]  ( .D(n538), .CPN(Clk_r), .Q(\Queue[3][30] ) );
  FDN1QM1P \Queue_reg[2][30]  ( .D(n506), .CPN(Clk_r), .Q(\Queue[2][30] ) );
  FDN1QM1P \Queue_reg[4][29]  ( .D(n409), .CPN(Clk_r), .Q(\Queue[4][29] ) );
  FDN1QM1P \Queue_reg[3][29]  ( .D(n537), .CPN(Clk_r), .Q(\Queue[3][29] ) );
  FDN1QM1P \Queue_reg[2][29]  ( .D(n505), .CPN(Clk_r), .Q(\Queue[2][29] ) );
  FDN1QM1P \Queue_reg[4][28]  ( .D(n408), .CPN(Clk_r), .Q(\Queue[4][28] ) );
  FDN1QM1P \Queue_reg[3][28]  ( .D(n536), .CPN(Clk_r), .Q(\Queue[3][28] ) );
  FDN1QM1P \Queue_reg[2][28]  ( .D(n504), .CPN(Clk_r), .Q(\Queue[2][28] ) );
  FDN1QM1P \Queue_reg[4][27]  ( .D(n407), .CPN(Clk_r), .Q(\Queue[4][27] ) );
  FDN1QM1P \Queue_reg[3][27]  ( .D(n535), .CPN(Clk_r), .Q(\Queue[3][27] ) );
  FDN1QM1P \Queue_reg[2][27]  ( .D(n503), .CPN(Clk_r), .Q(\Queue[2][27] ) );
  FDN1QM1P \Queue_reg[4][26]  ( .D(n406), .CPN(Clk_r), .Q(\Queue[4][26] ) );
  FDN1QM1P \Queue_reg[3][26]  ( .D(n534), .CPN(Clk_r), .Q(\Queue[3][26] ) );
  FDN1QM1P \Queue_reg[2][26]  ( .D(n502), .CPN(Clk_r), .Q(\Queue[2][26] ) );
  FDN1QM1P \Queue_reg[4][25]  ( .D(n405), .CPN(Clk_r), .Q(\Queue[4][25] ) );
  FDN1QM1P \Queue_reg[3][25]  ( .D(n533), .CPN(Clk_r), .Q(\Queue[3][25] ) );
  FDN1QM1P \Queue_reg[2][25]  ( .D(n501), .CPN(Clk_r), .Q(\Queue[2][25] ) );
  FDN1QM1P \Queue_reg[4][24]  ( .D(n404), .CPN(Clk_r), .Q(\Queue[4][24] ) );
  FDN1QM1P \Queue_reg[3][24]  ( .D(n532), .CPN(Clk_r), .Q(\Queue[3][24] ) );
  FDN1QM1P \Queue_reg[2][24]  ( .D(n500), .CPN(Clk_r), .Q(\Queue[2][24] ) );
  FDN1QM1P \Queue_reg[4][23]  ( .D(n403), .CPN(Clk_r), .Q(\Queue[4][23] ) );
  FDN1QM1P \Queue_reg[3][23]  ( .D(n531), .CPN(Clk_r), .Q(\Queue[3][23] ) );
  FDN1QM1P \Queue_reg[2][23]  ( .D(n499), .CPN(Clk_r), .Q(\Queue[2][23] ) );
  FDN1QM1P \Queue_reg[4][22]  ( .D(n402), .CPN(Clk_r), .Q(\Queue[4][22] ) );
  FDN1QM1P \Queue_reg[3][22]  ( .D(n530), .CPN(Clk_r), .Q(\Queue[3][22] ) );
  FDN1QM1P \Queue_reg[2][22]  ( .D(n498), .CPN(Clk_r), .Q(\Queue[2][22] ) );
  FDN1QM1P \Queue_reg[4][21]  ( .D(n401), .CPN(Clk_r), .Q(\Queue[4][21] ) );
  FDN1QM1P \Queue_reg[3][21]  ( .D(n529), .CPN(Clk_r), .Q(\Queue[3][21] ) );
  FDN1QM1P \Queue_reg[2][21]  ( .D(n497), .CPN(Clk_r), .Q(\Queue[2][21] ) );
  FDN1QM1P \Queue_reg[4][20]  ( .D(n400), .CPN(Clk_r), .Q(\Queue[4][20] ) );
  FDN1QM1P \Queue_reg[3][20]  ( .D(n528), .CPN(Clk_r), .Q(\Queue[3][20] ) );
  FDN1QM1P \Queue_reg[2][20]  ( .D(n496), .CPN(Clk_r), .Q(\Queue[2][20] ) );
  FDN1QM1P \Queue_reg[4][19]  ( .D(n399), .CPN(Clk_r), .Q(\Queue[4][19] ) );
  FDN1QM1P \Queue_reg[3][19]  ( .D(n527), .CPN(Clk_r), .Q(\Queue[3][19] ) );
  FDN1QM1P \Queue_reg[2][19]  ( .D(n495), .CPN(Clk_r), .Q(\Queue[2][19] ) );
  FDN1QM1P \Queue_reg[4][18]  ( .D(n398), .CPN(Clk_r), .Q(\Queue[4][18] ) );
  FDN1QM1P \Queue_reg[3][18]  ( .D(n526), .CPN(Clk_r), .Q(\Queue[3][18] ) );
  FDN1QM1P \Queue_reg[2][18]  ( .D(n494), .CPN(Clk_r), .Q(\Queue[2][18] ) );
  FDN1QM1P \Queue_reg[4][17]  ( .D(n397), .CPN(Clk_r), .Q(\Queue[4][17] ) );
  FDN1QM1P \Queue_reg[3][17]  ( .D(n525), .CPN(Clk_r), .Q(\Queue[3][17] ) );
  FDN1QM1P \Queue_reg[2][17]  ( .D(n493), .CPN(Clk_r), .Q(\Queue[2][17] ) );
  FDN1QM1P \Queue_reg[4][16]  ( .D(n396), .CPN(Clk_r), .Q(\Queue[4][16] ) );
  FDN1QM1P \Queue_reg[3][16]  ( .D(n524), .CPN(Clk_r), .Q(\Queue[3][16] ) );
  FDN1QM1P \Queue_reg[2][16]  ( .D(n492), .CPN(Clk_r), .Q(\Queue[2][16] ) );
  FDN1QM1P \Queue_reg[4][15]  ( .D(n395), .CPN(Clk_r), .Q(\Queue[4][15] ) );
  FDN1QM1P \Queue_reg[3][15]  ( .D(n523), .CPN(Clk_r), .Q(\Queue[3][15] ) );
  FDN1QM1P \Queue_reg[2][15]  ( .D(n491), .CPN(Clk_r), .Q(\Queue[2][15] ) );
  FDN1QM1P \Queue_reg[4][14]  ( .D(n394), .CPN(Clk_r), .Q(\Queue[4][14] ) );
  FDN1QM1P \Queue_reg[3][14]  ( .D(n522), .CPN(Clk_r), .Q(\Queue[3][14] ) );
  FDN1QM1P \Queue_reg[2][14]  ( .D(n490), .CPN(Clk_r), .Q(\Queue[2][14] ) );
  FDN1QM1P \Queue_reg[4][13]  ( .D(n393), .CPN(Clk_r), .Q(\Queue[4][13] ) );
  FDN1QM1P \Queue_reg[3][13]  ( .D(n521), .CPN(Clk_r), .Q(\Queue[3][13] ) );
  FDN1QM1P \Queue_reg[2][13]  ( .D(n489), .CPN(Clk_r), .Q(\Queue[2][13] ) );
  FDN1QM1P \Queue_reg[4][12]  ( .D(n392), .CPN(Clk_r), .Q(\Queue[4][12] ) );
  FDN1QM1P \Queue_reg[3][12]  ( .D(n520), .CPN(Clk_r), .Q(\Queue[3][12] ) );
  FDN1QM1P \Queue_reg[2][12]  ( .D(n488), .CPN(Clk_r), .Q(\Queue[2][12] ) );
  FDN1QM1P \Queue_reg[4][11]  ( .D(n391), .CPN(Clk_r), .Q(\Queue[4][11] ) );
  FDN1QM1P \Queue_reg[3][11]  ( .D(n519), .CPN(Clk_r), .Q(\Queue[3][11] ) );
  FDN1QM1P \Queue_reg[2][11]  ( .D(n487), .CPN(Clk_r), .Q(\Queue[2][11] ) );
  FDN1QM1P \Queue_reg[4][10]  ( .D(n390), .CPN(Clk_r), .Q(\Queue[4][10] ) );
  FDN1QM1P \Queue_reg[3][10]  ( .D(n518), .CPN(Clk_r), .Q(\Queue[3][10] ) );
  FDN1QM1P \Queue_reg[2][10]  ( .D(n486), .CPN(Clk_r), .Q(\Queue[2][10] ) );
  FDN1QM1P \Queue_reg[4][9]  ( .D(n389), .CPN(Clk_r), .Q(\Queue[4][9] ) );
  FDN1QM1P \Queue_reg[3][9]  ( .D(n517), .CPN(Clk_r), .Q(\Queue[3][9] ) );
  FDN1QM1P \Queue_reg[2][9]  ( .D(n485), .CPN(Clk_r), .Q(\Queue[2][9] ) );
  FDN1QM1P \Queue_reg[4][8]  ( .D(n388), .CPN(Clk_r), .Q(\Queue[4][8] ) );
  FDN1QM1P \Queue_reg[3][8]  ( .D(n516), .CPN(Clk_r), .Q(\Queue[3][8] ) );
  FDN1QM1P \Queue_reg[2][8]  ( .D(n484), .CPN(Clk_r), .Q(\Queue[2][8] ) );
  FDN1QM1P \Queue_reg[4][7]  ( .D(n387), .CPN(Clk_r), .Q(\Queue[4][7] ) );
  FDN1QM1P \Queue_reg[3][7]  ( .D(n515), .CPN(Clk_r), .Q(\Queue[3][7] ) );
  FDN1QM1P \Queue_reg[2][7]  ( .D(n483), .CPN(Clk_r), .Q(\Queue[2][7] ) );
  FDN1QM1P \Queue_reg[4][6]  ( .D(n386), .CPN(Clk_r), .Q(\Queue[4][6] ) );
  FDN1QM1P \Queue_reg[3][6]  ( .D(n514), .CPN(Clk_r), .Q(\Queue[3][6] ) );
  FDN1QM1P \Queue_reg[2][6]  ( .D(n482), .CPN(Clk_r), .Q(\Queue[2][6] ) );
  FDN1QM1P \Queue_reg[4][5]  ( .D(n385), .CPN(Clk_r), .Q(\Queue[4][5] ) );
  FDN1QM1P \Queue_reg[3][5]  ( .D(n513), .CPN(Clk_r), .Q(\Queue[3][5] ) );
  FDN1QM1P \Queue_reg[2][5]  ( .D(n481), .CPN(Clk_r), .Q(\Queue[2][5] ) );
  FDN1QM1P \Queue_reg[4][4]  ( .D(n384), .CPN(Clk_r), .Q(\Queue[4][4] ) );
  FDN1QM1P \Queue_reg[3][4]  ( .D(n512), .CPN(Clk_r), .Q(\Queue[3][4] ) );
  FDN1QM1P \Queue_reg[2][4]  ( .D(n480), .CPN(Clk_r), .Q(\Queue[2][4] ) );
  FDN1QM1P \Queue_reg[4][3]  ( .D(n383), .CPN(Clk_r), .Q(\Queue[4][3] ) );
  FDN1QM1P \Queue_reg[3][3]  ( .D(n511), .CPN(Clk_r), .Q(\Queue[3][3] ) );
  FDN1QM1P \Queue_reg[2][3]  ( .D(n479), .CPN(Clk_r), .Q(\Queue[2][3] ) );
  FDN1QM1P \Queue_reg[4][2]  ( .D(n382), .CPN(Clk_r), .Q(\Queue[4][2] ) );
  FDN1QM1P \Queue_reg[3][2]  ( .D(n510), .CPN(Clk_r), .Q(\Queue[3][2] ) );
  FDN1QM1P \Queue_reg[2][2]  ( .D(n478), .CPN(Clk_r), .Q(\Queue[2][2] ) );
  FDN1QM1P \Queue_reg[4][1]  ( .D(n381), .CPN(Clk_r), .Q(\Queue[4][1] ) );
  FDN1QM1P \Queue_reg[3][1]  ( .D(n509), .CPN(Clk_r), .Q(\Queue[3][1] ) );
  FDN1QM1P \Queue_reg[2][1]  ( .D(n477), .CPN(Clk_r), .Q(\Queue[2][1] ) );
  FDN1QM1P \Queue_reg[4][0]  ( .D(n380), .CPN(Clk_r), .Q(\Queue[4][0] ) );
  FDN1QM1P \Queue_reg[3][0]  ( .D(n508), .CPN(Clk_r), .Q(\Queue[3][0] ) );
  FDN1QM1P \Queue_reg[2][0]  ( .D(n476), .CPN(Clk_r), .Q(\Queue[2][0] ) );
  FDN1QM1P \Queue_reg[4][31]  ( .D(n379), .CPN(Clk_r), .Q(\Queue[4][31] ) );
  FDN1QM1P \Queue_reg[3][31]  ( .D(n539), .CPN(Clk_r), .Q(\Queue[3][31] ) );
  FDN1QM1P \Queue_reg[2][31]  ( .D(n507), .CPN(Clk_r), .Q(\Queue[2][31] ) );
  FDN2QM1P Full_reg ( .D(n411), .CPN(Clk_r), .CD(Rst_n), .Q(Full) );
  FDN1QM1P \Queue_reg[1][31]  ( .D(n443), .CPN(Clk_r), .Q(\Queue[1][31] ) );
  FDN1QM1P \Queue_reg[0][31]  ( .D(n475), .CPN(Clk_r), .Q(Packet_Out[31]) );
  FDN1QM1P \Queue_reg[1][30]  ( .D(n442), .CPN(Clk_r), .Q(\Queue[1][30] ) );
  FDN1QM1P \Queue_reg[0][30]  ( .D(n474), .CPN(Clk_r), .Q(Packet_Out[30]) );
  FDN1QM1P \Queue_reg[1][29]  ( .D(n441), .CPN(Clk_r), .Q(\Queue[1][29] ) );
  FDN1QM1P \Queue_reg[0][29]  ( .D(n473), .CPN(Clk_r), .Q(Packet_Out[29]) );
  FDN1QM1P \Queue_reg[1][28]  ( .D(n440), .CPN(Clk_r), .Q(\Queue[1][28] ) );
  FDN1QM1P \Queue_reg[0][28]  ( .D(n472), .CPN(Clk_r), .Q(Packet_Out[28]) );
  FDN1QM1P \Queue_reg[1][27]  ( .D(n439), .CPN(Clk_r), .Q(\Queue[1][27] ) );
  FDN1QM1P \Queue_reg[0][27]  ( .D(n471), .CPN(Clk_r), .Q(Packet_Out[27]) );
  FDN1QM1P \Queue_reg[1][26]  ( .D(n438), .CPN(Clk_r), .Q(\Queue[1][26] ) );
  FDN1QM1P \Queue_reg[0][26]  ( .D(n470), .CPN(Clk_r), .Q(Packet_Out[26]) );
  FDN1QM1P \Queue_reg[1][25]  ( .D(n437), .CPN(Clk_r), .Q(\Queue[1][25] ) );
  FDN1QM1P \Queue_reg[0][25]  ( .D(n469), .CPN(Clk_r), .Q(Packet_Out[25]) );
  FDN1QM1P \Queue_reg[1][24]  ( .D(n436), .CPN(Clk_r), .Q(\Queue[1][24] ) );
  FDN1QM1P \Queue_reg[0][24]  ( .D(n468), .CPN(Clk_r), .Q(Packet_Out[24]) );
  FDN1QM1P \Queue_reg[1][23]  ( .D(n435), .CPN(Clk_r), .Q(\Queue[1][23] ) );
  FDN1QM1P \Queue_reg[0][23]  ( .D(n467), .CPN(Clk_r), .Q(Packet_Out[23]) );
  FDN1QM1P \Queue_reg[1][22]  ( .D(n434), .CPN(Clk_r), .Q(\Queue[1][22] ) );
  FDN1QM1P \Queue_reg[0][22]  ( .D(n466), .CPN(Clk_r), .Q(Packet_Out[22]) );
  FDN1QM1P \Queue_reg[1][21]  ( .D(n433), .CPN(Clk_r), .Q(\Queue[1][21] ) );
  FDN1QM1P \Queue_reg[0][21]  ( .D(n465), .CPN(Clk_r), .Q(Packet_Out[21]) );
  FDN1QM1P \Queue_reg[1][20]  ( .D(n432), .CPN(Clk_r), .Q(\Queue[1][20] ) );
  FDN1QM1P \Queue_reg[0][20]  ( .D(n464), .CPN(Clk_r), .Q(Packet_Out[20]) );
  FDN1QM1P \Queue_reg[1][19]  ( .D(n431), .CPN(Clk_r), .Q(\Queue[1][19] ) );
  FDN1QM1P \Queue_reg[0][19]  ( .D(n463), .CPN(Clk_r), .Q(Packet_Out[19]) );
  FDN1QM1P \Queue_reg[1][18]  ( .D(n430), .CPN(Clk_r), .Q(\Queue[1][18] ) );
  FDN1QM1P \Queue_reg[0][18]  ( .D(n462), .CPN(Clk_r), .Q(Packet_Out[18]) );
  FDN1QM1P \Queue_reg[1][17]  ( .D(n429), .CPN(Clk_r), .Q(\Queue[1][17] ) );
  FDN1QM1P \Queue_reg[0][17]  ( .D(n461), .CPN(Clk_r), .Q(Packet_Out[17]) );
  FDN1QM1P \Queue_reg[1][16]  ( .D(n428), .CPN(Clk_r), .Q(\Queue[1][16] ) );
  FDN1QM1P \Queue_reg[0][16]  ( .D(n460), .CPN(Clk_r), .Q(Packet_Out[16]) );
  FDN1QM1P \Queue_reg[1][15]  ( .D(n427), .CPN(Clk_r), .Q(\Queue[1][15] ) );
  FDN1QM1P \Queue_reg[0][15]  ( .D(n459), .CPN(Clk_r), .Q(Packet_Out[15]) );
  FDN1QM1P \Queue_reg[1][14]  ( .D(n426), .CPN(Clk_r), .Q(\Queue[1][14] ) );
  FDN1QM1P \Queue_reg[0][14]  ( .D(n458), .CPN(Clk_r), .Q(Packet_Out[14]) );
  FDN1QM1P \Queue_reg[1][13]  ( .D(n425), .CPN(Clk_r), .Q(\Queue[1][13] ) );
  FDN1QM1P \Queue_reg[0][13]  ( .D(n457), .CPN(Clk_r), .Q(Packet_Out[13]) );
  FDN1QM1P \Queue_reg[1][12]  ( .D(n424), .CPN(Clk_r), .Q(\Queue[1][12] ) );
  FDN1QM1P \Queue_reg[0][12]  ( .D(n456), .CPN(Clk_r), .Q(Packet_Out[12]) );
  FDN1QM1P \Queue_reg[1][11]  ( .D(n423), .CPN(Clk_r), .Q(\Queue[1][11] ) );
  FDN1QM1P \Queue_reg[0][11]  ( .D(n455), .CPN(Clk_r), .Q(Packet_Out[11]) );
  FDN1QM1P \Queue_reg[1][10]  ( .D(n422), .CPN(Clk_r), .Q(\Queue[1][10] ) );
  FDN1QM1P \Queue_reg[0][10]  ( .D(n454), .CPN(Clk_r), .Q(Packet_Out[10]) );
  FDN1QM1P \Queue_reg[1][9]  ( .D(n421), .CPN(Clk_r), .Q(\Queue[1][9] ) );
  FDN1QM1P \Queue_reg[0][9]  ( .D(n453), .CPN(Clk_r), .Q(Packet_Out[9]) );
  FDN1QM1P \Queue_reg[1][8]  ( .D(n420), .CPN(Clk_r), .Q(\Queue[1][8] ) );
  FDN1QM1P \Queue_reg[0][8]  ( .D(n452), .CPN(Clk_r), .Q(Packet_Out[8]) );
  FDN1QM1P \Queue_reg[1][7]  ( .D(n419), .CPN(Clk_r), .Q(\Queue[1][7] ) );
  FDN1QM1P \Queue_reg[0][7]  ( .D(n451), .CPN(Clk_r), .Q(Packet_Out[7]) );
  FDN1QM1P \Queue_reg[1][6]  ( .D(n418), .CPN(Clk_r), .Q(\Queue[1][6] ) );
  FDN1QM1P \Queue_reg[0][6]  ( .D(n450), .CPN(Clk_r), .Q(Packet_Out[6]) );
  FDN1QM1P \Queue_reg[1][5]  ( .D(n417), .CPN(Clk_r), .Q(\Queue[1][5] ) );
  FDN1QM1P \Queue_reg[0][5]  ( .D(n449), .CPN(Clk_r), .Q(Packet_Out[5]) );
  FDN1QM1P \Queue_reg[1][4]  ( .D(n416), .CPN(Clk_r), .Q(\Queue[1][4] ) );
  FDN1QM1P \Queue_reg[0][4]  ( .D(n448), .CPN(Clk_r), .Q(Packet_Out[4]) );
  FDN1QM1P \Queue_reg[1][3]  ( .D(n415), .CPN(Clk_r), .Q(\Queue[1][3] ) );
  FDN1QM1P \Queue_reg[0][3]  ( .D(n447), .CPN(Clk_r), .Q(Packet_Out[3]) );
  FDN1QM1P \Queue_reg[1][2]  ( .D(n414), .CPN(Clk_r), .Q(\Queue[1][2] ) );
  FDN1QM1P \Queue_reg[0][2]  ( .D(n446), .CPN(Clk_r), .Q(Packet_Out[2]) );
  FDN1QM1P \Queue_reg[1][1]  ( .D(n413), .CPN(Clk_r), .Q(\Queue[1][1] ) );
  FDN1QM1P \Queue_reg[0][1]  ( .D(n445), .CPN(Clk_r), .Q(Packet_Out[1]) );
  FDN1QM1P \Queue_reg[1][0]  ( .D(n412), .CPN(Clk_r), .Q(\Queue[1][0] ) );
  FDN1QM1P \Queue_reg[0][0]  ( .D(n444), .CPN(Clk_r), .Q(Packet_Out[0]) );
  FDN2QM1P Empty_reg ( .D(n541), .CPN(Clk_r), .CD(Rst_n), .Q(n540) );
  BUFM2P U3 ( .A(n96), .Z(n10) );
  BUFM1P U4 ( .A(n96), .Z(n11) );
  BUFM2P U5 ( .A(n56), .Z(n5) );
  BUFM2P U6 ( .A(n131), .Z(n4) );
  BUFM2P U7 ( .A(n204), .Z(n3) );
  N1M1P U8 ( .A(Read_Ack), .Z(n136) );
  NR3M1P U9 ( .A(Count[0]), .B(Count[2]), .C(n21), .Z(n99) );
  NR3M1P U10 ( .A(Count[2]), .B(n22), .C(n21), .Z(n139) );
  NR3M1P U11 ( .A(n22), .B(Count[2]), .C(Count[1]), .Z(n375) );
  BUFM2P U12 ( .A(n94), .Z(n9) );
  NR2FM3P U13 ( .A(n60), .B(n20), .Z(n19) );
  OAI211M4P U14 ( .A(n139), .B(n138), .C(Rst_n), .D(n137), .Z(n205) );
  OAI211M4P U15 ( .A(n139), .B(n136), .C(n6), .D(n97), .Z(n134) );
  OAI211M4P U16 ( .A(n141), .B(n136), .C(n6), .D(n135), .Z(n207) );
  OAI21M2P U17 ( .A(n6), .B(Read_Ack), .C(n23), .Z(n55) );
  N1M2P U18 ( .A(n6), .Z(n98) );
  NR3M1P U19 ( .A(Count[0]), .B(Count[1]), .C(n18), .Z(n141) );
  N1M1P U20 ( .A(Count[0]), .Z(n22) );
  N1M1P U21 ( .A(Count[2]), .Z(n18) );
  N1M1P U22 ( .A(Count[1]), .Z(n21) );
  ND2M2P U23 ( .A(Read_Ack), .B(Rst_n), .Z(n140) );
  NR2M3P U24 ( .A(Read_Ack), .B(n98), .Z(n17) );
  BUFM10P U25 ( .A(Write_Ack), .Z(n6) );
  ND2M1P U26 ( .A(n17), .B(Rst_n), .Z(n60) );
  OAI211M4P U27 ( .A(n99), .B(n138), .C(Rst_n), .D(n137), .Z(n132) );
  N1M1P U28 ( .A(Packet_In[29]), .Z(n201) );
  N1M1P U29 ( .A(Packet_In[28]), .Z(n199) );
  N1M1P U30 ( .A(Packet_In[26]), .Z(n195) );
  N1M1P U31 ( .A(Packet_In[27]), .Z(n197) );
  N1M1P U32 ( .A(Packet_In[31]), .Z(n208) );
  N1M1P U33 ( .A(Packet_In[24]), .Z(n191) );
  N1M1P U34 ( .A(Packet_In[22]), .Z(n187) );
  N1M1P U35 ( .A(Packet_In[25]), .Z(n193) );
  N1M1P U36 ( .A(Packet_In[21]), .Z(n185) );
  N1M1P U37 ( .A(Packet_In[20]), .Z(n183) );
  N1M1P U38 ( .A(Packet_In[23]), .Z(n189) );
  N1M1P U39 ( .A(Packet_In[2]), .Z(n147) );
  N1M1P U40 ( .A(Packet_In[5]), .Z(n153) );
  N1M1P U41 ( .A(Packet_In[4]), .Z(n151) );
  N1M1P U42 ( .A(Packet_In[6]), .Z(n155) );
  N1M1P U43 ( .A(Packet_In[3]), .Z(n149) );
  N1M1P U44 ( .A(Packet_In[1]), .Z(n145) );
  N1M1P U45 ( .A(Packet_In[16]), .Z(n175) );
  N1M1P U46 ( .A(Packet_In[15]), .Z(n173) );
  N1M1P U47 ( .A(Packet_In[11]), .Z(n165) );
  N1M1P U48 ( .A(Packet_In[7]), .Z(n157) );
  N1M1P U49 ( .A(Packet_In[10]), .Z(n163) );
  N1M1P U50 ( .A(Packet_In[9]), .Z(n161) );
  N1M1P U51 ( .A(Packet_In[12]), .Z(n167) );
  N1M1P U52 ( .A(Packet_In[8]), .Z(n159) );
  N1M1P U53 ( .A(Packet_In[0]), .Z(n143) );
  N1M1P U54 ( .A(Packet_In[30]), .Z(n203) );
  N1M1P U55 ( .A(Packet_In[17]), .Z(n177) );
  N1M1P U56 ( .A(Packet_In[19]), .Z(n181) );
  N1M1P U57 ( .A(Packet_In[18]), .Z(n179) );
  N1M1P U58 ( .A(Packet_In[14]), .Z(n171) );
  N1M1P U59 ( .A(Packet_In[13]), .Z(n169) );
  BUFM2P U60 ( .A(n55), .Z(n7) );
  BUFM2P U61 ( .A(n55), .Z(n8) );
  N1M2P U62 ( .A(n61), .Z(n93) );
  OAI211M1P U63 ( .A(n375), .B(n136), .C(n6), .D(n61), .Z(n96) );
  N1M2P U64 ( .A(n17), .Z(n138) );
  OAI211M4P U65 ( .A(n99), .B(n136), .C(n6), .D(n23), .Z(n58) );
  NR2M1P U66 ( .A(n136), .B(n6), .Z(n374) );
  NR2M1P U67 ( .A(n17), .B(n374), .Z(n373) );
  AOI22CDNM1P U68 ( .A(n373), .B(n22), .C(n373), .D(n22), .Z(n376) );
  N1M1P U69 ( .A(n374), .Z(n16) );
  AOI22M1P U70 ( .A(Count[0]), .B(n138), .C(n16), .D(n22), .Z(n13) );
  AOI22CDNM1P U71 ( .A(Count[1]), .B(n13), .C(n13), .D(Count[1]), .Z(n377) );
  ND3M1P U72 ( .A(n22), .B(n18), .C(n21), .Z(n59) );
  ND2M1P U73 ( .A(Count[1]), .B(Read_Ack), .Z(n12) );
  OAI211M1P U74 ( .A(Count[1]), .B(n138), .C(n13), .D(n12), .Z(n14) );
  AOI22M1P U75 ( .A(n17), .B(n139), .C(Count[2]), .D(n14), .Z(n15) );
  OAI21M1P U76 ( .A(n59), .B(n16), .C(n15), .Z(n378) );
  N1M1P U77 ( .A(n141), .Z(n20) );
  AOI22CDNM1P U78 ( .A(n19), .B(n208), .C(\Queue[4][31] ), .D(n19), .Z(n379)
         );
  AOI22CDNM1P U79 ( .A(n19), .B(n143), .C(\Queue[4][0] ), .D(n19), .Z(n380) );
  AOI22CDNM1P U80 ( .A(n19), .B(n145), .C(\Queue[4][1] ), .D(n19), .Z(n381) );
  AOI22CDNM1P U81 ( .A(n19), .B(n147), .C(\Queue[4][2] ), .D(n19), .Z(n382) );
  AOI22CDNM1P U82 ( .A(n19), .B(n149), .C(\Queue[4][3] ), .D(n19), .Z(n383) );
  AOI22CDNM1P U83 ( .A(n19), .B(n151), .C(\Queue[4][4] ), .D(n19), .Z(n384) );
  AOI22CDNM1P U84 ( .A(n19), .B(n153), .C(\Queue[4][5] ), .D(n19), .Z(n385) );
  AOI22CDNM1P U85 ( .A(n19), .B(n155), .C(\Queue[4][6] ), .D(n19), .Z(n386) );
  AOI22CDNM1P U86 ( .A(n19), .B(n157), .C(\Queue[4][7] ), .D(n19), .Z(n387) );
  AOI22CDNM1P U87 ( .A(n19), .B(n159), .C(\Queue[4][8] ), .D(n19), .Z(n388) );
  AOI22CDNM1P U88 ( .A(n19), .B(n161), .C(\Queue[4][9] ), .D(n19), .Z(n389) );
  AOI22CDNM1P U89 ( .A(n19), .B(n163), .C(\Queue[4][10] ), .D(n19), .Z(n390)
         );
  AOI22CDNM1P U90 ( .A(n19), .B(n165), .C(\Queue[4][11] ), .D(n19), .Z(n391)
         );
  AOI22CDNM1P U91 ( .A(n19), .B(n167), .C(\Queue[4][12] ), .D(n19), .Z(n392)
         );
  AOI22CDNM1P U92 ( .A(n19), .B(n169), .C(\Queue[4][13] ), .D(n19), .Z(n393)
         );
  AOI22CDNM1P U93 ( .A(n19), .B(n171), .C(\Queue[4][14] ), .D(n19), .Z(n394)
         );
  AOI22CDNM1P U94 ( .A(n19), .B(n173), .C(\Queue[4][15] ), .D(n19), .Z(n395)
         );
  AOI22CDNM1P U95 ( .A(n19), .B(n175), .C(\Queue[4][16] ), .D(n19), .Z(n396)
         );
  AOI22CDNM1P U96 ( .A(n19), .B(n177), .C(\Queue[4][17] ), .D(n19), .Z(n397)
         );
  AOI22CDNM1P U97 ( .A(n19), .B(n179), .C(\Queue[4][18] ), .D(n19), .Z(n398)
         );
  AOI22CDNM1P U98 ( .A(n19), .B(n181), .C(\Queue[4][19] ), .D(n19), .Z(n399)
         );
  AOI22CDNM1P U99 ( .A(n19), .B(n183), .C(\Queue[4][20] ), .D(n19), .Z(n400)
         );
  AOI22CDNM1P U100 ( .A(n19), .B(n185), .C(\Queue[4][21] ), .D(n19), .Z(n401)
         );
  AOI22CDNM1P U101 ( .A(n19), .B(n187), .C(\Queue[4][22] ), .D(n19), .Z(n402)
         );
  AOI22CDNM1P U102 ( .A(n19), .B(n189), .C(\Queue[4][23] ), .D(n19), .Z(n403)
         );
  AOI22CDNM1P U103 ( .A(n19), .B(n191), .C(\Queue[4][24] ), .D(n19), .Z(n404)
         );
  AOI22CDNM1P U104 ( .A(n19), .B(n193), .C(\Queue[4][25] ), .D(n19), .Z(n405)
         );
  AOI22CDNM1P U105 ( .A(n19), .B(n195), .C(\Queue[4][26] ), .D(n19), .Z(n406)
         );
  AOI22CDNM1P U106 ( .A(n19), .B(n197), .C(\Queue[4][27] ), .D(n19), .Z(n407)
         );
  AOI22CDNM1P U107 ( .A(n19), .B(n199), .C(\Queue[4][28] ), .D(n19), .Z(n408)
         );
  AOI22CDNM1P U108 ( .A(n19), .B(n201), .C(\Queue[4][29] ), .D(n19), .Z(n409)
         );
  AOI22CDNM1P U109 ( .A(n19), .B(n203), .C(\Queue[4][30] ), .D(n19), .Z(n410)
         );
  OAI22CDNM1P U110 ( .A(n138), .B(n20), .C(n373), .D(Full), .Z(n411) );
  OA21M1P U111 ( .A(n138), .B(n375), .C(Rst_n), .Z(n23) );
  AOI21M1P U112 ( .A(n6), .B(n99), .C(n140), .Z(n56) );
  AOI22M1P U113 ( .A(\Queue[2][0] ), .B(n5), .C(\Queue[1][0] ), .D(n7), .Z(n24) );
  OAI21M1P U114 ( .A(n143), .B(n58), .C(n24), .Z(n412) );
  AOI22M1P U115 ( .A(n5), .B(\Queue[2][1] ), .C(\Queue[1][1] ), .D(n7), .Z(n25) );
  OAI21M1P U116 ( .A(n58), .B(n145), .C(n25), .Z(n413) );
  AOI22M1P U117 ( .A(n5), .B(\Queue[2][2] ), .C(\Queue[1][2] ), .D(n7), .Z(n26) );
  OAI21M1P U118 ( .A(n58), .B(n147), .C(n26), .Z(n414) );
  AOI22M1P U119 ( .A(n5), .B(\Queue[2][3] ), .C(\Queue[1][3] ), .D(n7), .Z(n27) );
  OAI21M1P U120 ( .A(n58), .B(n149), .C(n27), .Z(n415) );
  AOI22M1P U121 ( .A(n5), .B(\Queue[2][4] ), .C(\Queue[1][4] ), .D(n7), .Z(n28) );
  OAI21M1P U122 ( .A(n58), .B(n151), .C(n28), .Z(n416) );
  AOI22M1P U123 ( .A(n5), .B(\Queue[2][5] ), .C(\Queue[1][5] ), .D(n7), .Z(n29) );
  OAI21M1P U124 ( .A(n58), .B(n153), .C(n29), .Z(n417) );
  AOI22M1P U125 ( .A(n5), .B(\Queue[2][6] ), .C(\Queue[1][6] ), .D(n7), .Z(n30) );
  OAI21M1P U126 ( .A(n58), .B(n155), .C(n30), .Z(n418) );
  AOI22M1P U127 ( .A(n5), .B(\Queue[2][7] ), .C(\Queue[1][7] ), .D(n7), .Z(n31) );
  OAI21M1P U128 ( .A(n58), .B(n157), .C(n31), .Z(n419) );
  AOI22M1P U129 ( .A(n5), .B(\Queue[2][8] ), .C(\Queue[1][8] ), .D(n7), .Z(n32) );
  OAI21M1P U130 ( .A(n58), .B(n159), .C(n32), .Z(n420) );
  AOI22M1P U131 ( .A(n5), .B(\Queue[2][9] ), .C(\Queue[1][9] ), .D(n55), .Z(
        n33) );
  OAI21M1P U132 ( .A(n58), .B(n161), .C(n33), .Z(n421) );
  AOI22M1P U133 ( .A(n5), .B(\Queue[2][10] ), .C(\Queue[1][10] ), .D(n55), .Z(
        n34) );
  OAI21M1P U134 ( .A(n58), .B(n163), .C(n34), .Z(n422) );
  AOI22M1P U135 ( .A(n5), .B(\Queue[2][11] ), .C(\Queue[1][11] ), .D(n55), .Z(
        n35) );
  OAI21M1P U136 ( .A(n58), .B(n165), .C(n35), .Z(n423) );
  AOI22M1P U137 ( .A(n5), .B(\Queue[2][12] ), .C(\Queue[1][12] ), .D(n55), .Z(
        n36) );
  OAI21M1P U138 ( .A(n58), .B(n167), .C(n36), .Z(n424) );
  AOI22M1P U139 ( .A(n5), .B(\Queue[2][13] ), .C(\Queue[1][13] ), .D(n55), .Z(
        n37) );
  OAI21M1P U140 ( .A(n58), .B(n169), .C(n37), .Z(n425) );
  AOI22M1P U141 ( .A(n5), .B(\Queue[2][14] ), .C(\Queue[1][14] ), .D(n55), .Z(
        n38) );
  OAI21M1P U142 ( .A(n58), .B(n171), .C(n38), .Z(n426) );
  AOI22M1P U143 ( .A(n5), .B(\Queue[2][15] ), .C(\Queue[1][15] ), .D(n8), .Z(
        n39) );
  OAI21M1P U144 ( .A(n58), .B(n173), .C(n39), .Z(n427) );
  AOI22M1P U145 ( .A(n5), .B(\Queue[2][16] ), .C(\Queue[1][16] ), .D(n7), .Z(
        n40) );
  OAI21M1P U146 ( .A(n58), .B(n175), .C(n40), .Z(n428) );
  AOI22M1P U147 ( .A(n5), .B(\Queue[2][17] ), .C(\Queue[1][17] ), .D(n8), .Z(
        n41) );
  OAI21M1P U148 ( .A(n58), .B(n177), .C(n41), .Z(n429) );
  AOI22M1P U149 ( .A(n5), .B(\Queue[2][18] ), .C(\Queue[1][18] ), .D(n8), .Z(
        n42) );
  OAI21M1P U150 ( .A(n58), .B(n179), .C(n42), .Z(n430) );
  AOI22M1P U151 ( .A(n5), .B(\Queue[2][19] ), .C(\Queue[1][19] ), .D(n8), .Z(
        n43) );
  OAI21M1P U152 ( .A(n58), .B(n181), .C(n43), .Z(n431) );
  AOI22M1P U153 ( .A(n5), .B(\Queue[2][20] ), .C(\Queue[1][20] ), .D(n8), .Z(
        n44) );
  OAI21M1P U154 ( .A(n58), .B(n183), .C(n44), .Z(n432) );
  AOI22M1P U155 ( .A(n5), .B(\Queue[2][21] ), .C(\Queue[1][21] ), .D(n8), .Z(
        n45) );
  OAI21M1P U156 ( .A(n58), .B(n185), .C(n45), .Z(n433) );
  AOI22M1P U157 ( .A(n5), .B(\Queue[2][22] ), .C(\Queue[1][22] ), .D(n8), .Z(
        n46) );
  OAI21M1P U158 ( .A(n58), .B(n187), .C(n46), .Z(n434) );
  AOI22M1P U159 ( .A(n5), .B(\Queue[2][23] ), .C(\Queue[1][23] ), .D(n8), .Z(
        n47) );
  OAI21M1P U160 ( .A(n58), .B(n189), .C(n47), .Z(n435) );
  AOI22M1P U161 ( .A(n5), .B(\Queue[2][24] ), .C(\Queue[1][24] ), .D(n8), .Z(
        n48) );
  OAI21M1P U162 ( .A(n58), .B(n191), .C(n48), .Z(n436) );
  AOI22M1P U163 ( .A(n5), .B(\Queue[2][25] ), .C(\Queue[1][25] ), .D(n8), .Z(
        n49) );
  OAI21M1P U164 ( .A(n58), .B(n193), .C(n49), .Z(n437) );
  AOI22M1P U165 ( .A(n5), .B(\Queue[2][26] ), .C(\Queue[1][26] ), .D(n8), .Z(
        n50) );
  OAI21M1P U166 ( .A(n58), .B(n195), .C(n50), .Z(n438) );
  AOI22M1P U167 ( .A(n5), .B(\Queue[2][27] ), .C(\Queue[1][27] ), .D(n8), .Z(
        n51) );
  OAI21M1P U168 ( .A(n58), .B(n197), .C(n51), .Z(n439) );
  AOI22M1P U169 ( .A(n5), .B(\Queue[2][28] ), .C(\Queue[1][28] ), .D(n7), .Z(
        n52) );
  OAI21M1P U170 ( .A(n58), .B(n199), .C(n52), .Z(n440) );
  AOI22M1P U171 ( .A(n5), .B(\Queue[2][29] ), .C(\Queue[1][29] ), .D(n55), .Z(
        n53) );
  OAI21M1P U172 ( .A(n58), .B(n201), .C(n53), .Z(n441) );
  AOI22M1P U173 ( .A(n5), .B(\Queue[2][30] ), .C(\Queue[1][30] ), .D(n8), .Z(
        n54) );
  OAI21M1P U174 ( .A(n58), .B(n203), .C(n54), .Z(n442) );
  AOI22M1P U175 ( .A(n5), .B(\Queue[2][31] ), .C(\Queue[1][31] ), .D(n7), .Z(
        n57) );
  OAI21M1P U176 ( .A(n58), .B(n208), .C(n57), .Z(n443) );
  OAI21M1P U177 ( .A(n60), .B(n59), .C(n140), .Z(n61) );
  AOI21M1P U178 ( .A(n6), .B(n375), .C(n140), .Z(n94) );
  AOI22M1P U179 ( .A(\Queue[1][0] ), .B(n94), .C(n93), .D(Packet_Out[0]), .Z(
        n62) );
  OAI21M1P U180 ( .A(n143), .B(n10), .C(n62), .Z(n444) );
  AOI22M1P U181 ( .A(\Queue[1][1] ), .B(n94), .C(n93), .D(Packet_Out[1]), .Z(
        n63) );
  OAI21M1P U182 ( .A(n145), .B(n10), .C(n63), .Z(n445) );
  AOI22M1P U183 ( .A(\Queue[1][2] ), .B(n94), .C(n93), .D(Packet_Out[2]), .Z(
        n64) );
  OAI21M1P U184 ( .A(n147), .B(n10), .C(n64), .Z(n446) );
  AOI22M1P U185 ( .A(\Queue[1][3] ), .B(n94), .C(n93), .D(Packet_Out[3]), .Z(
        n65) );
  OAI21M1P U186 ( .A(n149), .B(n10), .C(n65), .Z(n447) );
  AOI22M1P U187 ( .A(\Queue[1][4] ), .B(n94), .C(n93), .D(Packet_Out[4]), .Z(
        n66) );
  OAI21M1P U188 ( .A(n151), .B(n10), .C(n66), .Z(n448) );
  AOI22M1P U189 ( .A(\Queue[1][5] ), .B(n94), .C(n93), .D(Packet_Out[5]), .Z(
        n67) );
  OAI21M1P U190 ( .A(n153), .B(n10), .C(n67), .Z(n449) );
  AOI22M1P U191 ( .A(\Queue[1][6] ), .B(n9), .C(n93), .D(Packet_Out[6]), .Z(
        n68) );
  OAI21M1P U192 ( .A(n155), .B(n10), .C(n68), .Z(n450) );
  AOI22M1P U193 ( .A(\Queue[1][7] ), .B(n9), .C(n93), .D(Packet_Out[7]), .Z(
        n69) );
  OAI21M1P U194 ( .A(n157), .B(n10), .C(n69), .Z(n451) );
  AOI22M1P U195 ( .A(\Queue[1][8] ), .B(n9), .C(n93), .D(Packet_Out[8]), .Z(
        n70) );
  OAI21M1P U196 ( .A(n159), .B(n10), .C(n70), .Z(n452) );
  AOI22M1P U197 ( .A(\Queue[1][9] ), .B(n9), .C(n93), .D(Packet_Out[9]), .Z(
        n71) );
  OAI21M1P U198 ( .A(n161), .B(n10), .C(n71), .Z(n453) );
  AOI22M1P U199 ( .A(\Queue[1][10] ), .B(n9), .C(n93), .D(Packet_Out[10]), .Z(
        n72) );
  OAI21M1P U200 ( .A(n163), .B(n10), .C(n72), .Z(n454) );
  AOI22M1P U201 ( .A(\Queue[1][11] ), .B(n9), .C(n93), .D(Packet_Out[11]), .Z(
        n73) );
  OAI21M1P U202 ( .A(n165), .B(n10), .C(n73), .Z(n455) );
  AOI22M1P U203 ( .A(\Queue[1][12] ), .B(n9), .C(n93), .D(Packet_Out[12]), .Z(
        n74) );
  OAI21M1P U204 ( .A(n167), .B(n10), .C(n74), .Z(n456) );
  AOI22M1P U205 ( .A(\Queue[1][13] ), .B(n9), .C(n93), .D(Packet_Out[13]), .Z(
        n75) );
  OAI21M1P U206 ( .A(n169), .B(n10), .C(n75), .Z(n457) );
  AOI22M1P U207 ( .A(\Queue[1][14] ), .B(n9), .C(n93), .D(Packet_Out[14]), .Z(
        n76) );
  OAI21M1P U208 ( .A(n171), .B(n10), .C(n76), .Z(n458) );
  AOI22M1P U209 ( .A(\Queue[1][15] ), .B(n9), .C(n93), .D(Packet_Out[15]), .Z(
        n77) );
  OAI21M1P U210 ( .A(n173), .B(n10), .C(n77), .Z(n459) );
  AOI22M1P U211 ( .A(\Queue[1][16] ), .B(n9), .C(n93), .D(Packet_Out[16]), .Z(
        n78) );
  OAI21M1P U212 ( .A(n175), .B(n10), .C(n78), .Z(n460) );
  AOI22M1P U213 ( .A(\Queue[1][17] ), .B(n9), .C(n93), .D(Packet_Out[17]), .Z(
        n79) );
  OAI21M1P U214 ( .A(n177), .B(n10), .C(n79), .Z(n461) );
  AOI22M1P U215 ( .A(\Queue[1][18] ), .B(n9), .C(n93), .D(Packet_Out[18]), .Z(
        n80) );
  OAI21M1P U216 ( .A(n179), .B(n10), .C(n80), .Z(n462) );
  AOI22M1P U217 ( .A(\Queue[1][19] ), .B(n9), .C(n93), .D(Packet_Out[19]), .Z(
        n81) );
  OAI21M1P U218 ( .A(n181), .B(n10), .C(n81), .Z(n463) );
  AOI22M1P U219 ( .A(\Queue[1][20] ), .B(n9), .C(n93), .D(Packet_Out[20]), .Z(
        n82) );
  OAI21M1P U220 ( .A(n183), .B(n11), .C(n82), .Z(n464) );
  AOI22M1P U221 ( .A(\Queue[1][21] ), .B(n9), .C(n93), .D(Packet_Out[21]), .Z(
        n83) );
  OAI21M1P U222 ( .A(n185), .B(n11), .C(n83), .Z(n465) );
  AOI22M1P U223 ( .A(\Queue[1][22] ), .B(n9), .C(n93), .D(Packet_Out[22]), .Z(
        n84) );
  OAI21M1P U224 ( .A(n187), .B(n11), .C(n84), .Z(n466) );
  AOI22M1P U225 ( .A(\Queue[1][23] ), .B(n9), .C(n93), .D(Packet_Out[23]), .Z(
        n85) );
  OAI21M1P U226 ( .A(n189), .B(n11), .C(n85), .Z(n467) );
  AOI22M1P U227 ( .A(\Queue[1][24] ), .B(n9), .C(n93), .D(Packet_Out[24]), .Z(
        n86) );
  OAI21M1P U228 ( .A(n191), .B(n11), .C(n86), .Z(n468) );
  AOI22M1P U229 ( .A(\Queue[1][25] ), .B(n9), .C(n93), .D(Packet_Out[25]), .Z(
        n87) );
  OAI21M1P U230 ( .A(n193), .B(n11), .C(n87), .Z(n469) );
  AOI22M1P U231 ( .A(\Queue[1][26] ), .B(n9), .C(n93), .D(Packet_Out[26]), .Z(
        n88) );
  OAI21M1P U232 ( .A(n195), .B(n11), .C(n88), .Z(n470) );
  AOI22M1P U233 ( .A(\Queue[1][27] ), .B(n9), .C(n93), .D(Packet_Out[27]), .Z(
        n89) );
  OAI21M1P U234 ( .A(n197), .B(n11), .C(n89), .Z(n471) );
  AOI22M1P U235 ( .A(\Queue[1][28] ), .B(n9), .C(n93), .D(Packet_Out[28]), .Z(
        n90) );
  OAI21M1P U236 ( .A(n199), .B(n11), .C(n90), .Z(n472) );
  AOI22M1P U237 ( .A(\Queue[1][29] ), .B(n9), .C(n93), .D(Packet_Out[29]), .Z(
        n91) );
  OAI21M1P U238 ( .A(n201), .B(n11), .C(n91), .Z(n473) );
  AOI22M1P U239 ( .A(\Queue[1][30] ), .B(n9), .C(n93), .D(Packet_Out[30]), .Z(
        n92) );
  OAI21M1P U240 ( .A(n203), .B(n10), .C(n92), .Z(n474) );
  AOI22M1P U241 ( .A(\Queue[1][31] ), .B(n9), .C(n93), .D(Packet_Out[31]), .Z(
        n95) );
  OAI21M1P U242 ( .A(n208), .B(n11), .C(n95), .Z(n475) );
  OA21M1P U243 ( .A(n138), .B(n99), .C(Rst_n), .Z(n97) );
  ND2M1P U244 ( .A(n98), .B(n136), .Z(n137) );
  AOI21M1P U245 ( .A(n6), .B(n139), .C(n140), .Z(n131) );
  AOI22M1P U246 ( .A(\Queue[2][0] ), .B(n132), .C(\Queue[3][0] ), .D(n4), .Z(
        n100) );
  OAI21M1P U247 ( .A(n143), .B(n134), .C(n100), .Z(n476) );
  AOI22M1P U248 ( .A(\Queue[2][1] ), .B(n132), .C(n4), .D(\Queue[3][1] ), .Z(
        n101) );
  OAI21M1P U249 ( .A(n145), .B(n134), .C(n101), .Z(n477) );
  AOI22M1P U250 ( .A(\Queue[2][2] ), .B(n132), .C(n4), .D(\Queue[3][2] ), .Z(
        n102) );
  OAI21M1P U251 ( .A(n147), .B(n134), .C(n102), .Z(n478) );
  AOI22M1P U252 ( .A(\Queue[2][3] ), .B(n132), .C(n4), .D(\Queue[3][3] ), .Z(
        n103) );
  OAI21M1P U253 ( .A(n149), .B(n134), .C(n103), .Z(n479) );
  AOI22M1P U254 ( .A(\Queue[2][4] ), .B(n132), .C(n4), .D(\Queue[3][4] ), .Z(
        n104) );
  OAI21M1P U255 ( .A(n151), .B(n134), .C(n104), .Z(n480) );
  AOI22M1P U256 ( .A(\Queue[2][5] ), .B(n132), .C(n4), .D(\Queue[3][5] ), .Z(
        n105) );
  OAI21M1P U257 ( .A(n153), .B(n134), .C(n105), .Z(n481) );
  AOI22M1P U258 ( .A(\Queue[2][6] ), .B(n132), .C(n4), .D(\Queue[3][6] ), .Z(
        n106) );
  OAI21M1P U259 ( .A(n155), .B(n134), .C(n106), .Z(n482) );
  AOI22M1P U260 ( .A(\Queue[2][7] ), .B(n132), .C(n4), .D(\Queue[3][7] ), .Z(
        n107) );
  OAI21M1P U261 ( .A(n157), .B(n134), .C(n107), .Z(n483) );
  AOI22M1P U262 ( .A(\Queue[2][8] ), .B(n132), .C(n4), .D(\Queue[3][8] ), .Z(
        n108) );
  OAI21M1P U263 ( .A(n159), .B(n134), .C(n108), .Z(n484) );
  AOI22M1P U264 ( .A(\Queue[2][9] ), .B(n132), .C(n4), .D(\Queue[3][9] ), .Z(
        n109) );
  OAI21M1P U265 ( .A(n161), .B(n134), .C(n109), .Z(n485) );
  AOI22M1P U266 ( .A(\Queue[2][10] ), .B(n132), .C(n4), .D(\Queue[3][10] ), 
        .Z(n110) );
  OAI21M1P U267 ( .A(n163), .B(n134), .C(n110), .Z(n486) );
  AOI22M1P U268 ( .A(\Queue[2][11] ), .B(n132), .C(n4), .D(\Queue[3][11] ), 
        .Z(n111) );
  OAI21M1P U269 ( .A(n165), .B(n134), .C(n111), .Z(n487) );
  AOI22M1P U270 ( .A(\Queue[2][12] ), .B(n132), .C(n4), .D(\Queue[3][12] ), 
        .Z(n112) );
  OAI21M1P U271 ( .A(n167), .B(n134), .C(n112), .Z(n488) );
  AOI22M1P U272 ( .A(\Queue[2][13] ), .B(n132), .C(n4), .D(\Queue[3][13] ), 
        .Z(n113) );
  OAI21M1P U273 ( .A(n169), .B(n134), .C(n113), .Z(n489) );
  AOI22M1P U274 ( .A(\Queue[2][14] ), .B(n132), .C(n4), .D(\Queue[3][14] ), 
        .Z(n114) );
  OAI21M1P U275 ( .A(n171), .B(n134), .C(n114), .Z(n490) );
  AOI22M1P U276 ( .A(\Queue[2][15] ), .B(n132), .C(n4), .D(\Queue[3][15] ), 
        .Z(n115) );
  OAI21M1P U277 ( .A(n173), .B(n134), .C(n115), .Z(n491) );
  AOI22M1P U278 ( .A(\Queue[2][16] ), .B(n132), .C(n4), .D(\Queue[3][16] ), 
        .Z(n116) );
  OAI21M1P U279 ( .A(n175), .B(n134), .C(n116), .Z(n492) );
  AOI22M1P U280 ( .A(\Queue[2][17] ), .B(n132), .C(n4), .D(\Queue[3][17] ), 
        .Z(n117) );
  OAI21M1P U281 ( .A(n177), .B(n134), .C(n117), .Z(n493) );
  AOI22M1P U282 ( .A(\Queue[2][18] ), .B(n132), .C(n4), .D(\Queue[3][18] ), 
        .Z(n118) );
  OAI21M1P U283 ( .A(n179), .B(n134), .C(n118), .Z(n494) );
  AOI22M1P U284 ( .A(\Queue[2][19] ), .B(n132), .C(n4), .D(\Queue[3][19] ), 
        .Z(n119) );
  OAI21M1P U285 ( .A(n181), .B(n134), .C(n119), .Z(n495) );
  AOI22M1P U286 ( .A(\Queue[2][20] ), .B(n132), .C(n4), .D(\Queue[3][20] ), 
        .Z(n120) );
  OAI21M1P U287 ( .A(n183), .B(n134), .C(n120), .Z(n496) );
  AOI22M1P U288 ( .A(\Queue[2][21] ), .B(n132), .C(n4), .D(\Queue[3][21] ), 
        .Z(n121) );
  OAI21M1P U289 ( .A(n185), .B(n134), .C(n121), .Z(n497) );
  AOI22M1P U290 ( .A(\Queue[2][22] ), .B(n132), .C(n4), .D(\Queue[3][22] ), 
        .Z(n122) );
  OAI21M1P U291 ( .A(n187), .B(n134), .C(n122), .Z(n498) );
  AOI22M1P U292 ( .A(\Queue[2][23] ), .B(n132), .C(n4), .D(\Queue[3][23] ), 
        .Z(n123) );
  OAI21M1P U293 ( .A(n189), .B(n134), .C(n123), .Z(n499) );
  AOI22M1P U294 ( .A(\Queue[2][24] ), .B(n132), .C(n4), .D(\Queue[3][24] ), 
        .Z(n124) );
  OAI21M1P U295 ( .A(n191), .B(n134), .C(n124), .Z(n500) );
  AOI22M1P U296 ( .A(\Queue[2][25] ), .B(n132), .C(n4), .D(\Queue[3][25] ), 
        .Z(n125) );
  OAI21M1P U297 ( .A(n193), .B(n134), .C(n125), .Z(n501) );
  AOI22M1P U298 ( .A(\Queue[2][26] ), .B(n132), .C(n4), .D(\Queue[3][26] ), 
        .Z(n126) );
  OAI21M1P U299 ( .A(n195), .B(n134), .C(n126), .Z(n502) );
  AOI22M1P U300 ( .A(\Queue[2][27] ), .B(n132), .C(n4), .D(\Queue[3][27] ), 
        .Z(n127) );
  OAI21M1P U301 ( .A(n197), .B(n134), .C(n127), .Z(n503) );
  AOI22M1P U302 ( .A(\Queue[2][28] ), .B(n132), .C(n4), .D(\Queue[3][28] ), 
        .Z(n128) );
  OAI21M1P U303 ( .A(n199), .B(n134), .C(n128), .Z(n504) );
  AOI22M1P U304 ( .A(\Queue[2][29] ), .B(n132), .C(n4), .D(\Queue[3][29] ), 
        .Z(n129) );
  OAI21M1P U305 ( .A(n201), .B(n134), .C(n129), .Z(n505) );
  AOI22M1P U306 ( .A(\Queue[2][30] ), .B(n132), .C(n4), .D(\Queue[3][30] ), 
        .Z(n130) );
  OAI21M1P U307 ( .A(n203), .B(n134), .C(n130), .Z(n506) );
  AOI22M1P U308 ( .A(\Queue[2][31] ), .B(n132), .C(n4), .D(\Queue[3][31] ), 
        .Z(n133) );
  OAI21M1P U309 ( .A(n208), .B(n134), .C(n133), .Z(n507) );
  OA21M1P U310 ( .A(n138), .B(n139), .C(Rst_n), .Z(n135) );
  AOI21M1P U311 ( .A(n6), .B(n141), .C(n140), .Z(n204) );
  AOI22M1P U312 ( .A(\Queue[3][0] ), .B(n205), .C(n3), .D(\Queue[4][0] ), .Z(
        n142) );
  OAI21M1P U313 ( .A(n143), .B(n207), .C(n142), .Z(n508) );
  AOI22M1P U314 ( .A(\Queue[3][1] ), .B(n205), .C(n3), .D(\Queue[4][1] ), .Z(
        n144) );
  OAI21M1P U315 ( .A(n145), .B(n207), .C(n144), .Z(n509) );
  AOI22M1P U316 ( .A(\Queue[3][2] ), .B(n205), .C(n3), .D(\Queue[4][2] ), .Z(
        n146) );
  OAI21M1P U317 ( .A(n147), .B(n207), .C(n146), .Z(n510) );
  AOI22M1P U318 ( .A(\Queue[3][3] ), .B(n205), .C(n3), .D(\Queue[4][3] ), .Z(
        n148) );
  OAI21M1P U319 ( .A(n149), .B(n207), .C(n148), .Z(n511) );
  AOI22M1P U320 ( .A(\Queue[3][4] ), .B(n205), .C(n3), .D(\Queue[4][4] ), .Z(
        n150) );
  OAI21M1P U321 ( .A(n151), .B(n207), .C(n150), .Z(n512) );
  AOI22M1P U322 ( .A(\Queue[3][5] ), .B(n205), .C(n3), .D(\Queue[4][5] ), .Z(
        n152) );
  OAI21M1P U323 ( .A(n153), .B(n207), .C(n152), .Z(n513) );
  AOI22M1P U324 ( .A(\Queue[3][6] ), .B(n205), .C(n3), .D(\Queue[4][6] ), .Z(
        n154) );
  OAI21M1P U325 ( .A(n155), .B(n207), .C(n154), .Z(n514) );
  AOI22M1P U326 ( .A(\Queue[3][7] ), .B(n205), .C(n3), .D(\Queue[4][7] ), .Z(
        n156) );
  OAI21M1P U327 ( .A(n157), .B(n207), .C(n156), .Z(n515) );
  AOI22M1P U328 ( .A(\Queue[3][8] ), .B(n205), .C(n3), .D(\Queue[4][8] ), .Z(
        n158) );
  OAI21M1P U329 ( .A(n159), .B(n207), .C(n158), .Z(n516) );
  AOI22M1P U330 ( .A(\Queue[3][9] ), .B(n205), .C(n3), .D(\Queue[4][9] ), .Z(
        n160) );
  OAI21M1P U331 ( .A(n161), .B(n207), .C(n160), .Z(n517) );
  AOI22M1P U332 ( .A(\Queue[3][10] ), .B(n205), .C(n3), .D(\Queue[4][10] ), 
        .Z(n162) );
  OAI21M1P U333 ( .A(n163), .B(n207), .C(n162), .Z(n518) );
  AOI22M1P U334 ( .A(\Queue[3][11] ), .B(n205), .C(n3), .D(\Queue[4][11] ), 
        .Z(n164) );
  OAI21M1P U335 ( .A(n165), .B(n207), .C(n164), .Z(n519) );
  AOI22M1P U336 ( .A(\Queue[3][12] ), .B(n205), .C(n3), .D(\Queue[4][12] ), 
        .Z(n166) );
  OAI21M1P U337 ( .A(n167), .B(n207), .C(n166), .Z(n520) );
  AOI22M1P U338 ( .A(\Queue[3][13] ), .B(n205), .C(n3), .D(\Queue[4][13] ), 
        .Z(n168) );
  OAI21M1P U339 ( .A(n169), .B(n207), .C(n168), .Z(n521) );
  AOI22M1P U340 ( .A(\Queue[3][14] ), .B(n205), .C(n3), .D(\Queue[4][14] ), 
        .Z(n170) );
  OAI21M1P U341 ( .A(n171), .B(n207), .C(n170), .Z(n522) );
  AOI22M1P U342 ( .A(\Queue[3][15] ), .B(n205), .C(n3), .D(\Queue[4][15] ), 
        .Z(n172) );
  OAI21M1P U343 ( .A(n173), .B(n207), .C(n172), .Z(n523) );
  AOI22M1P U344 ( .A(\Queue[3][16] ), .B(n205), .C(n3), .D(\Queue[4][16] ), 
        .Z(n174) );
  OAI21M1P U345 ( .A(n175), .B(n207), .C(n174), .Z(n524) );
  AOI22M1P U346 ( .A(\Queue[3][17] ), .B(n205), .C(n3), .D(\Queue[4][17] ), 
        .Z(n176) );
  OAI21M1P U347 ( .A(n177), .B(n207), .C(n176), .Z(n525) );
  AOI22M1P U348 ( .A(\Queue[3][18] ), .B(n205), .C(n3), .D(\Queue[4][18] ), 
        .Z(n178) );
  OAI21M1P U349 ( .A(n179), .B(n207), .C(n178), .Z(n526) );
  AOI22M1P U350 ( .A(\Queue[3][19] ), .B(n205), .C(n3), .D(\Queue[4][19] ), 
        .Z(n180) );
  OAI21M1P U351 ( .A(n181), .B(n207), .C(n180), .Z(n527) );
  AOI22M1P U352 ( .A(\Queue[3][20] ), .B(n205), .C(n3), .D(\Queue[4][20] ), 
        .Z(n182) );
  OAI21M1P U353 ( .A(n183), .B(n207), .C(n182), .Z(n528) );
  AOI22M1P U354 ( .A(\Queue[3][21] ), .B(n205), .C(n3), .D(\Queue[4][21] ), 
        .Z(n184) );
  OAI21M1P U355 ( .A(n185), .B(n207), .C(n184), .Z(n529) );
  AOI22M1P U356 ( .A(\Queue[3][22] ), .B(n205), .C(n3), .D(\Queue[4][22] ), 
        .Z(n186) );
  OAI21M1P U357 ( .A(n187), .B(n207), .C(n186), .Z(n530) );
  AOI22M1P U358 ( .A(\Queue[3][23] ), .B(n205), .C(n3), .D(\Queue[4][23] ), 
        .Z(n188) );
  OAI21M1P U359 ( .A(n189), .B(n207), .C(n188), .Z(n531) );
  AOI22M1P U360 ( .A(\Queue[3][24] ), .B(n205), .C(n3), .D(\Queue[4][24] ), 
        .Z(n190) );
  OAI21M1P U361 ( .A(n191), .B(n207), .C(n190), .Z(n532) );
  AOI22M1P U362 ( .A(\Queue[3][25] ), .B(n205), .C(n3), .D(\Queue[4][25] ), 
        .Z(n192) );
  OAI21M1P U363 ( .A(n193), .B(n207), .C(n192), .Z(n533) );
  AOI22M1P U364 ( .A(\Queue[3][26] ), .B(n205), .C(n3), .D(\Queue[4][26] ), 
        .Z(n194) );
  OAI21M1P U365 ( .A(n195), .B(n207), .C(n194), .Z(n534) );
  AOI22M1P U366 ( .A(\Queue[3][27] ), .B(n205), .C(n3), .D(\Queue[4][27] ), 
        .Z(n196) );
  OAI21M1P U367 ( .A(n197), .B(n207), .C(n196), .Z(n535) );
  AOI22M1P U368 ( .A(\Queue[3][28] ), .B(n205), .C(n3), .D(\Queue[4][28] ), 
        .Z(n198) );
  OAI21M1P U369 ( .A(n199), .B(n207), .C(n198), .Z(n536) );
  AOI22M1P U370 ( .A(\Queue[3][29] ), .B(n205), .C(n3), .D(\Queue[4][29] ), 
        .Z(n200) );
  OAI21M1P U371 ( .A(n201), .B(n207), .C(n200), .Z(n537) );
  AOI22M1P U372 ( .A(\Queue[3][30] ), .B(n205), .C(n3), .D(\Queue[4][30] ), 
        .Z(n202) );
  OAI21M1P U373 ( .A(n203), .B(n207), .C(n202), .Z(n538) );
  AOI22M1P U374 ( .A(\Queue[3][31] ), .B(n205), .C(n3), .D(\Queue[4][31] ), 
        .Z(n206) );
  OAI21M1P U375 ( .A(n208), .B(n207), .C(n206), .Z(n539) );
  N1M1P U376 ( .A(n540), .Z(Empty) );
  AOI22M1P U377 ( .A(n375), .B(n374), .C(n373), .D(Empty), .Z(n541) );
endmodule


module Link_Control_1 ( Clk_r, Rst_n, Tx_Ready, Tx_Error, RxData_Valid, RxData, 
        Packet_From_Core, TxQueue_Write, RxQueue_Read, TxData_Valid, TxData, 
        Error_Ack, Core_Rcv_Ready, Packet_To_Core, RxQueue_Empty, TxQueue_Full
 );
  input [31:0] RxData;
  input [31:0] Packet_From_Core;
  output [31:0] TxData;
  output [31:0] Packet_To_Core;
  input Clk_r, Rst_n, Tx_Ready, Tx_Error, RxData_Valid, TxQueue_Write,
         RxQueue_Read;
  output TxData_Valid, Error_Ack, Core_Rcv_Ready, RxQueue_Empty, TxQueue_Full;
  wire   TxQueue_Read, TxQueue_Empty, RxQueue_Write, RxQueue_Full, N9, N16, n5,
         n6, n7, n8, n9;

  Packet_Queue_4 TxQueue ( .Clk_r(Clk_r), .Rst_n(Rst_n), .Packet_In(
        Packet_From_Core), .Read_Ack(TxQueue_Read), .Write_Ack(TxQueue_Write), 
        .Packet_Out(TxData), .Empty(TxQueue_Empty), .Full(TxQueue_Full) );
  Packet_Queue_3 RxQueue ( .Clk_r(Clk_r), .Rst_n(Rst_n), .Packet_In(RxData), 
        .Read_Ack(RxQueue_Read), .Write_Ack(RxQueue_Write), .Packet_Out(
        Packet_To_Core), .Empty(RxQueue_Empty), .Full(RxQueue_Full) );
  FD2QM1P Core_Rcv_Ready_reg ( .D(N9), .CP(Clk_r), .CD(Rst_n), .Q(
        Core_Rcv_Ready) );
  FD2QM1P TxQueue_Read_reg ( .D(N16), .CP(Clk_r), .CD(Rst_n), .Q(TxQueue_Read)
         );
  FD2QM1P Error_Ack_reg ( .D(Tx_Error), .CP(Clk_r), .CD(Rst_n), .Q(Error_Ack)
         );
  FD4QM1P RxQueue_Write_reg ( .D(n7), .CP(Clk_r), .SD(Rst_n), .Q(n6) );
  FD4QM1P TxData_Valid_reg ( .D(n9), .CP(Clk_r), .SD(Rst_n), .Q(n8) );
  N1M2P U3 ( .A(n6), .Z(RxQueue_Write) );
  NR2M1P U4 ( .A(n8), .B(Tx_Ready), .Z(N16) );
  NR2M1P U5 ( .A(RxData_Valid), .B(RxQueue_Full), .Z(n5) );
  OA21M1P U6 ( .A(Core_Rcv_Ready), .B(n5), .C(n6), .Z(N9) );
  N1M1P U7 ( .A(n8), .Z(TxData_Valid) );
  ND3M1P U8 ( .A(n6), .B(Core_Rcv_Ready), .C(RxData_Valid), .Z(n7) );
  AO21CNM1P U9 ( .A(n8), .B(TxQueue_Empty), .C(Tx_Ready), .Z(n9) );
endmodule


module Packet_Queue_5 ( Clk_r, Rst_n, Packet_In, Read_Ack, Write_Ack, 
        Packet_Out, Empty, Full );
  input [31:0] Packet_In;
  output [31:0] Packet_Out;
  input Clk_r, Rst_n, Read_Ack, Write_Ack;
  output Empty, Full;
  wire   \Queue[4][31] , \Queue[4][30] , \Queue[4][29] , \Queue[4][28] ,
         \Queue[4][27] , \Queue[4][26] , \Queue[4][25] , \Queue[4][24] ,
         \Queue[4][23] , \Queue[4][22] , \Queue[4][21] , \Queue[4][20] ,
         \Queue[4][19] , \Queue[4][18] , \Queue[4][17] , \Queue[4][16] ,
         \Queue[4][15] , \Queue[4][14] , \Queue[4][13] , \Queue[4][12] ,
         \Queue[4][11] , \Queue[4][10] , \Queue[4][9] , \Queue[4][8] ,
         \Queue[4][7] , \Queue[4][6] , \Queue[4][5] , \Queue[4][4] ,
         \Queue[4][3] , \Queue[4][2] , \Queue[4][1] , \Queue[4][0] ,
         \Queue[3][31] , \Queue[3][30] , \Queue[3][29] , \Queue[3][28] ,
         \Queue[3][27] , \Queue[3][26] , \Queue[3][25] , \Queue[3][24] ,
         \Queue[3][23] , \Queue[3][22] , \Queue[3][21] , \Queue[3][20] ,
         \Queue[3][19] , \Queue[3][18] , \Queue[3][17] , \Queue[3][16] ,
         \Queue[3][15] , \Queue[3][14] , \Queue[3][13] , \Queue[3][12] ,
         \Queue[3][11] , \Queue[3][10] , \Queue[3][9] , \Queue[3][8] ,
         \Queue[3][7] , \Queue[3][6] , \Queue[3][5] , \Queue[3][4] ,
         \Queue[3][3] , \Queue[3][2] , \Queue[3][1] , \Queue[3][0] ,
         \Queue[2][31] , \Queue[2][30] , \Queue[2][29] , \Queue[2][28] ,
         \Queue[2][27] , \Queue[2][26] , \Queue[2][25] , \Queue[2][24] ,
         \Queue[2][23] , \Queue[2][22] , \Queue[2][21] , \Queue[2][20] ,
         \Queue[2][19] , \Queue[2][18] , \Queue[2][17] , \Queue[2][16] ,
         \Queue[2][15] , \Queue[2][14] , \Queue[2][13] , \Queue[2][12] ,
         \Queue[2][11] , \Queue[2][10] , \Queue[2][9] , \Queue[2][8] ,
         \Queue[2][7] , \Queue[2][6] , \Queue[2][5] , \Queue[2][4] ,
         \Queue[2][3] , \Queue[2][2] , \Queue[2][1] , \Queue[2][0] ,
         \Queue[1][31] , \Queue[1][30] , \Queue[1][29] , \Queue[1][28] ,
         \Queue[1][27] , \Queue[1][26] , \Queue[1][25] , \Queue[1][24] ,
         \Queue[1][23] , \Queue[1][22] , \Queue[1][21] , \Queue[1][20] ,
         \Queue[1][19] , \Queue[1][18] , \Queue[1][17] , \Queue[1][16] ,
         \Queue[1][15] , \Queue[1][14] , \Queue[1][13] , \Queue[1][12] ,
         \Queue[1][11] , \Queue[1][10] , \Queue[1][9] , \Queue[1][8] ,
         \Queue[1][7] , \Queue[1][6] , \Queue[1][5] , \Queue[1][4] ,
         \Queue[1][3] , \Queue[1][2] , \Queue[1][1] , \Queue[1][0] , n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541;
  wire   [2:0] Count;

  FDN2QM1P \Count_reg[0]  ( .D(n376), .CPN(Clk_r), .CD(Rst_n), .Q(Count[0]) );
  FDN2QM1P \Count_reg[1]  ( .D(n377), .CPN(Clk_r), .CD(Rst_n), .Q(Count[1]) );
  FDN2QM1P \Count_reg[2]  ( .D(n378), .CPN(Clk_r), .CD(Rst_n), .Q(Count[2]) );
  FDN1QM1P \Queue_reg[4][30]  ( .D(n410), .CPN(Clk_r), .Q(\Queue[4][30] ) );
  FDN1QM1P \Queue_reg[3][30]  ( .D(n538), .CPN(Clk_r), .Q(\Queue[3][30] ) );
  FDN1QM1P \Queue_reg[2][30]  ( .D(n506), .CPN(Clk_r), .Q(\Queue[2][30] ) );
  FDN1QM1P \Queue_reg[4][29]  ( .D(n409), .CPN(Clk_r), .Q(\Queue[4][29] ) );
  FDN1QM1P \Queue_reg[3][29]  ( .D(n537), .CPN(Clk_r), .Q(\Queue[3][29] ) );
  FDN1QM1P \Queue_reg[2][29]  ( .D(n505), .CPN(Clk_r), .Q(\Queue[2][29] ) );
  FDN1QM1P \Queue_reg[4][28]  ( .D(n408), .CPN(Clk_r), .Q(\Queue[4][28] ) );
  FDN1QM1P \Queue_reg[3][28]  ( .D(n536), .CPN(Clk_r), .Q(\Queue[3][28] ) );
  FDN1QM1P \Queue_reg[2][28]  ( .D(n504), .CPN(Clk_r), .Q(\Queue[2][28] ) );
  FDN1QM1P \Queue_reg[4][27]  ( .D(n407), .CPN(Clk_r), .Q(\Queue[4][27] ) );
  FDN1QM1P \Queue_reg[3][27]  ( .D(n535), .CPN(Clk_r), .Q(\Queue[3][27] ) );
  FDN1QM1P \Queue_reg[2][27]  ( .D(n503), .CPN(Clk_r), .Q(\Queue[2][27] ) );
  FDN1QM1P \Queue_reg[4][26]  ( .D(n406), .CPN(Clk_r), .Q(\Queue[4][26] ) );
  FDN1QM1P \Queue_reg[3][26]  ( .D(n534), .CPN(Clk_r), .Q(\Queue[3][26] ) );
  FDN1QM1P \Queue_reg[2][26]  ( .D(n502), .CPN(Clk_r), .Q(\Queue[2][26] ) );
  FDN1QM1P \Queue_reg[4][25]  ( .D(n405), .CPN(Clk_r), .Q(\Queue[4][25] ) );
  FDN1QM1P \Queue_reg[3][25]  ( .D(n533), .CPN(Clk_r), .Q(\Queue[3][25] ) );
  FDN1QM1P \Queue_reg[2][25]  ( .D(n501), .CPN(Clk_r), .Q(\Queue[2][25] ) );
  FDN1QM1P \Queue_reg[4][24]  ( .D(n404), .CPN(Clk_r), .Q(\Queue[4][24] ) );
  FDN1QM1P \Queue_reg[3][24]  ( .D(n532), .CPN(Clk_r), .Q(\Queue[3][24] ) );
  FDN1QM1P \Queue_reg[2][24]  ( .D(n500), .CPN(Clk_r), .Q(\Queue[2][24] ) );
  FDN1QM1P \Queue_reg[4][23]  ( .D(n403), .CPN(Clk_r), .Q(\Queue[4][23] ) );
  FDN1QM1P \Queue_reg[3][23]  ( .D(n531), .CPN(Clk_r), .Q(\Queue[3][23] ) );
  FDN1QM1P \Queue_reg[2][23]  ( .D(n499), .CPN(Clk_r), .Q(\Queue[2][23] ) );
  FDN1QM1P \Queue_reg[4][22]  ( .D(n402), .CPN(Clk_r), .Q(\Queue[4][22] ) );
  FDN1QM1P \Queue_reg[3][22]  ( .D(n530), .CPN(Clk_r), .Q(\Queue[3][22] ) );
  FDN1QM1P \Queue_reg[2][22]  ( .D(n498), .CPN(Clk_r), .Q(\Queue[2][22] ) );
  FDN1QM1P \Queue_reg[4][21]  ( .D(n401), .CPN(Clk_r), .Q(\Queue[4][21] ) );
  FDN1QM1P \Queue_reg[3][21]  ( .D(n529), .CPN(Clk_r), .Q(\Queue[3][21] ) );
  FDN1QM1P \Queue_reg[2][21]  ( .D(n497), .CPN(Clk_r), .Q(\Queue[2][21] ) );
  FDN1QM1P \Queue_reg[4][20]  ( .D(n400), .CPN(Clk_r), .Q(\Queue[4][20] ) );
  FDN1QM1P \Queue_reg[3][20]  ( .D(n528), .CPN(Clk_r), .Q(\Queue[3][20] ) );
  FDN1QM1P \Queue_reg[2][20]  ( .D(n496), .CPN(Clk_r), .Q(\Queue[2][20] ) );
  FDN1QM1P \Queue_reg[4][19]  ( .D(n399), .CPN(Clk_r), .Q(\Queue[4][19] ) );
  FDN1QM1P \Queue_reg[3][19]  ( .D(n527), .CPN(Clk_r), .Q(\Queue[3][19] ) );
  FDN1QM1P \Queue_reg[2][19]  ( .D(n495), .CPN(Clk_r), .Q(\Queue[2][19] ) );
  FDN1QM1P \Queue_reg[4][18]  ( .D(n398), .CPN(Clk_r), .Q(\Queue[4][18] ) );
  FDN1QM1P \Queue_reg[3][18]  ( .D(n526), .CPN(Clk_r), .Q(\Queue[3][18] ) );
  FDN1QM1P \Queue_reg[2][18]  ( .D(n494), .CPN(Clk_r), .Q(\Queue[2][18] ) );
  FDN1QM1P \Queue_reg[4][17]  ( .D(n397), .CPN(Clk_r), .Q(\Queue[4][17] ) );
  FDN1QM1P \Queue_reg[3][17]  ( .D(n525), .CPN(Clk_r), .Q(\Queue[3][17] ) );
  FDN1QM1P \Queue_reg[2][17]  ( .D(n493), .CPN(Clk_r), .Q(\Queue[2][17] ) );
  FDN1QM1P \Queue_reg[4][16]  ( .D(n396), .CPN(Clk_r), .Q(\Queue[4][16] ) );
  FDN1QM1P \Queue_reg[3][16]  ( .D(n524), .CPN(Clk_r), .Q(\Queue[3][16] ) );
  FDN1QM1P \Queue_reg[2][16]  ( .D(n492), .CPN(Clk_r), .Q(\Queue[2][16] ) );
  FDN1QM1P \Queue_reg[4][15]  ( .D(n395), .CPN(Clk_r), .Q(\Queue[4][15] ) );
  FDN1QM1P \Queue_reg[3][15]  ( .D(n523), .CPN(Clk_r), .Q(\Queue[3][15] ) );
  FDN1QM1P \Queue_reg[2][15]  ( .D(n491), .CPN(Clk_r), .Q(\Queue[2][15] ) );
  FDN1QM1P \Queue_reg[4][14]  ( .D(n394), .CPN(Clk_r), .Q(\Queue[4][14] ) );
  FDN1QM1P \Queue_reg[3][14]  ( .D(n522), .CPN(Clk_r), .Q(\Queue[3][14] ) );
  FDN1QM1P \Queue_reg[2][14]  ( .D(n490), .CPN(Clk_r), .Q(\Queue[2][14] ) );
  FDN1QM1P \Queue_reg[4][13]  ( .D(n393), .CPN(Clk_r), .Q(\Queue[4][13] ) );
  FDN1QM1P \Queue_reg[3][13]  ( .D(n521), .CPN(Clk_r), .Q(\Queue[3][13] ) );
  FDN1QM1P \Queue_reg[2][13]  ( .D(n489), .CPN(Clk_r), .Q(\Queue[2][13] ) );
  FDN1QM1P \Queue_reg[4][12]  ( .D(n392), .CPN(Clk_r), .Q(\Queue[4][12] ) );
  FDN1QM1P \Queue_reg[3][12]  ( .D(n520), .CPN(Clk_r), .Q(\Queue[3][12] ) );
  FDN1QM1P \Queue_reg[2][12]  ( .D(n488), .CPN(Clk_r), .Q(\Queue[2][12] ) );
  FDN1QM1P \Queue_reg[4][11]  ( .D(n391), .CPN(Clk_r), .Q(\Queue[4][11] ) );
  FDN1QM1P \Queue_reg[3][11]  ( .D(n519), .CPN(Clk_r), .Q(\Queue[3][11] ) );
  FDN1QM1P \Queue_reg[2][11]  ( .D(n487), .CPN(Clk_r), .Q(\Queue[2][11] ) );
  FDN1QM1P \Queue_reg[4][10]  ( .D(n390), .CPN(Clk_r), .Q(\Queue[4][10] ) );
  FDN1QM1P \Queue_reg[3][10]  ( .D(n518), .CPN(Clk_r), .Q(\Queue[3][10] ) );
  FDN1QM1P \Queue_reg[2][10]  ( .D(n486), .CPN(Clk_r), .Q(\Queue[2][10] ) );
  FDN1QM1P \Queue_reg[4][9]  ( .D(n389), .CPN(Clk_r), .Q(\Queue[4][9] ) );
  FDN1QM1P \Queue_reg[3][9]  ( .D(n517), .CPN(Clk_r), .Q(\Queue[3][9] ) );
  FDN1QM1P \Queue_reg[2][9]  ( .D(n485), .CPN(Clk_r), .Q(\Queue[2][9] ) );
  FDN1QM1P \Queue_reg[4][8]  ( .D(n388), .CPN(Clk_r), .Q(\Queue[4][8] ) );
  FDN1QM1P \Queue_reg[3][8]  ( .D(n516), .CPN(Clk_r), .Q(\Queue[3][8] ) );
  FDN1QM1P \Queue_reg[2][8]  ( .D(n484), .CPN(Clk_r), .Q(\Queue[2][8] ) );
  FDN1QM1P \Queue_reg[4][7]  ( .D(n387), .CPN(Clk_r), .Q(\Queue[4][7] ) );
  FDN1QM1P \Queue_reg[3][7]  ( .D(n515), .CPN(Clk_r), .Q(\Queue[3][7] ) );
  FDN1QM1P \Queue_reg[2][7]  ( .D(n483), .CPN(Clk_r), .Q(\Queue[2][7] ) );
  FDN1QM1P \Queue_reg[4][6]  ( .D(n386), .CPN(Clk_r), .Q(\Queue[4][6] ) );
  FDN1QM1P \Queue_reg[3][6]  ( .D(n514), .CPN(Clk_r), .Q(\Queue[3][6] ) );
  FDN1QM1P \Queue_reg[2][6]  ( .D(n482), .CPN(Clk_r), .Q(\Queue[2][6] ) );
  FDN1QM1P \Queue_reg[4][5]  ( .D(n385), .CPN(Clk_r), .Q(\Queue[4][5] ) );
  FDN1QM1P \Queue_reg[3][5]  ( .D(n513), .CPN(Clk_r), .Q(\Queue[3][5] ) );
  FDN1QM1P \Queue_reg[2][5]  ( .D(n481), .CPN(Clk_r), .Q(\Queue[2][5] ) );
  FDN1QM1P \Queue_reg[4][4]  ( .D(n384), .CPN(Clk_r), .Q(\Queue[4][4] ) );
  FDN1QM1P \Queue_reg[3][4]  ( .D(n512), .CPN(Clk_r), .Q(\Queue[3][4] ) );
  FDN1QM1P \Queue_reg[2][4]  ( .D(n480), .CPN(Clk_r), .Q(\Queue[2][4] ) );
  FDN1QM1P \Queue_reg[4][3]  ( .D(n383), .CPN(Clk_r), .Q(\Queue[4][3] ) );
  FDN1QM1P \Queue_reg[3][3]  ( .D(n511), .CPN(Clk_r), .Q(\Queue[3][3] ) );
  FDN1QM1P \Queue_reg[2][3]  ( .D(n479), .CPN(Clk_r), .Q(\Queue[2][3] ) );
  FDN1QM1P \Queue_reg[4][2]  ( .D(n382), .CPN(Clk_r), .Q(\Queue[4][2] ) );
  FDN1QM1P \Queue_reg[3][2]  ( .D(n510), .CPN(Clk_r), .Q(\Queue[3][2] ) );
  FDN1QM1P \Queue_reg[2][2]  ( .D(n478), .CPN(Clk_r), .Q(\Queue[2][2] ) );
  FDN1QM1P \Queue_reg[4][1]  ( .D(n381), .CPN(Clk_r), .Q(\Queue[4][1] ) );
  FDN1QM1P \Queue_reg[3][1]  ( .D(n509), .CPN(Clk_r), .Q(\Queue[3][1] ) );
  FDN1QM1P \Queue_reg[2][1]  ( .D(n477), .CPN(Clk_r), .Q(\Queue[2][1] ) );
  FDN1QM1P \Queue_reg[4][0]  ( .D(n380), .CPN(Clk_r), .Q(\Queue[4][0] ) );
  FDN1QM1P \Queue_reg[3][0]  ( .D(n508), .CPN(Clk_r), .Q(\Queue[3][0] ) );
  FDN1QM1P \Queue_reg[2][0]  ( .D(n476), .CPN(Clk_r), .Q(\Queue[2][0] ) );
  FDN1QM1P \Queue_reg[4][31]  ( .D(n379), .CPN(Clk_r), .Q(\Queue[4][31] ) );
  FDN1QM1P \Queue_reg[3][31]  ( .D(n539), .CPN(Clk_r), .Q(\Queue[3][31] ) );
  FDN1QM1P \Queue_reg[2][31]  ( .D(n507), .CPN(Clk_r), .Q(\Queue[2][31] ) );
  FDN2QM1P Full_reg ( .D(n411), .CPN(Clk_r), .CD(Rst_n), .Q(Full) );
  FDN1QM1P \Queue_reg[1][31]  ( .D(n443), .CPN(Clk_r), .Q(\Queue[1][31] ) );
  FDN1QM1P \Queue_reg[0][31]  ( .D(n475), .CPN(Clk_r), .Q(Packet_Out[31]) );
  FDN1QM1P \Queue_reg[1][30]  ( .D(n442), .CPN(Clk_r), .Q(\Queue[1][30] ) );
  FDN1QM1P \Queue_reg[0][30]  ( .D(n474), .CPN(Clk_r), .Q(Packet_Out[30]) );
  FDN1QM1P \Queue_reg[1][29]  ( .D(n441), .CPN(Clk_r), .Q(\Queue[1][29] ) );
  FDN1QM1P \Queue_reg[0][29]  ( .D(n473), .CPN(Clk_r), .Q(Packet_Out[29]) );
  FDN1QM1P \Queue_reg[1][28]  ( .D(n440), .CPN(Clk_r), .Q(\Queue[1][28] ) );
  FDN1QM1P \Queue_reg[0][28]  ( .D(n472), .CPN(Clk_r), .Q(Packet_Out[28]) );
  FDN1QM1P \Queue_reg[1][27]  ( .D(n439), .CPN(Clk_r), .Q(\Queue[1][27] ) );
  FDN1QM1P \Queue_reg[0][27]  ( .D(n471), .CPN(Clk_r), .Q(Packet_Out[27]) );
  FDN1QM1P \Queue_reg[1][26]  ( .D(n438), .CPN(Clk_r), .Q(\Queue[1][26] ) );
  FDN1QM1P \Queue_reg[0][26]  ( .D(n470), .CPN(Clk_r), .Q(Packet_Out[26]) );
  FDN1QM1P \Queue_reg[1][25]  ( .D(n437), .CPN(Clk_r), .Q(\Queue[1][25] ) );
  FDN1QM1P \Queue_reg[0][25]  ( .D(n469), .CPN(Clk_r), .Q(Packet_Out[25]) );
  FDN1QM1P \Queue_reg[1][24]  ( .D(n436), .CPN(Clk_r), .Q(\Queue[1][24] ) );
  FDN1QM1P \Queue_reg[0][24]  ( .D(n468), .CPN(Clk_r), .Q(Packet_Out[24]) );
  FDN1QM1P \Queue_reg[1][23]  ( .D(n435), .CPN(Clk_r), .Q(\Queue[1][23] ) );
  FDN1QM1P \Queue_reg[0][23]  ( .D(n467), .CPN(Clk_r), .Q(Packet_Out[23]) );
  FDN1QM1P \Queue_reg[1][22]  ( .D(n434), .CPN(Clk_r), .Q(\Queue[1][22] ) );
  FDN1QM1P \Queue_reg[0][22]  ( .D(n466), .CPN(Clk_r), .Q(Packet_Out[22]) );
  FDN1QM1P \Queue_reg[1][21]  ( .D(n433), .CPN(Clk_r), .Q(\Queue[1][21] ) );
  FDN1QM1P \Queue_reg[0][21]  ( .D(n465), .CPN(Clk_r), .Q(Packet_Out[21]) );
  FDN1QM1P \Queue_reg[1][20]  ( .D(n432), .CPN(Clk_r), .Q(\Queue[1][20] ) );
  FDN1QM1P \Queue_reg[0][20]  ( .D(n464), .CPN(Clk_r), .Q(Packet_Out[20]) );
  FDN1QM1P \Queue_reg[1][19]  ( .D(n431), .CPN(Clk_r), .Q(\Queue[1][19] ) );
  FDN1QM1P \Queue_reg[0][19]  ( .D(n463), .CPN(Clk_r), .Q(Packet_Out[19]) );
  FDN1QM1P \Queue_reg[1][18]  ( .D(n430), .CPN(Clk_r), .Q(\Queue[1][18] ) );
  FDN1QM1P \Queue_reg[0][18]  ( .D(n462), .CPN(Clk_r), .Q(Packet_Out[18]) );
  FDN1QM1P \Queue_reg[1][17]  ( .D(n429), .CPN(Clk_r), .Q(\Queue[1][17] ) );
  FDN1QM1P \Queue_reg[0][17]  ( .D(n461), .CPN(Clk_r), .Q(Packet_Out[17]) );
  FDN1QM1P \Queue_reg[1][16]  ( .D(n428), .CPN(Clk_r), .Q(\Queue[1][16] ) );
  FDN1QM1P \Queue_reg[0][16]  ( .D(n460), .CPN(Clk_r), .Q(Packet_Out[16]) );
  FDN1QM1P \Queue_reg[1][15]  ( .D(n427), .CPN(Clk_r), .Q(\Queue[1][15] ) );
  FDN1QM1P \Queue_reg[0][15]  ( .D(n459), .CPN(Clk_r), .Q(Packet_Out[15]) );
  FDN1QM1P \Queue_reg[1][14]  ( .D(n426), .CPN(Clk_r), .Q(\Queue[1][14] ) );
  FDN1QM1P \Queue_reg[0][14]  ( .D(n458), .CPN(Clk_r), .Q(Packet_Out[14]) );
  FDN1QM1P \Queue_reg[1][13]  ( .D(n425), .CPN(Clk_r), .Q(\Queue[1][13] ) );
  FDN1QM1P \Queue_reg[0][13]  ( .D(n457), .CPN(Clk_r), .Q(Packet_Out[13]) );
  FDN1QM1P \Queue_reg[1][12]  ( .D(n424), .CPN(Clk_r), .Q(\Queue[1][12] ) );
  FDN1QM1P \Queue_reg[0][12]  ( .D(n456), .CPN(Clk_r), .Q(Packet_Out[12]) );
  FDN1QM1P \Queue_reg[1][11]  ( .D(n423), .CPN(Clk_r), .Q(\Queue[1][11] ) );
  FDN1QM1P \Queue_reg[0][11]  ( .D(n455), .CPN(Clk_r), .Q(Packet_Out[11]) );
  FDN1QM1P \Queue_reg[1][10]  ( .D(n422), .CPN(Clk_r), .Q(\Queue[1][10] ) );
  FDN1QM1P \Queue_reg[0][10]  ( .D(n454), .CPN(Clk_r), .Q(Packet_Out[10]) );
  FDN1QM1P \Queue_reg[1][9]  ( .D(n421), .CPN(Clk_r), .Q(\Queue[1][9] ) );
  FDN1QM1P \Queue_reg[0][9]  ( .D(n453), .CPN(Clk_r), .Q(Packet_Out[9]) );
  FDN1QM1P \Queue_reg[1][8]  ( .D(n420), .CPN(Clk_r), .Q(\Queue[1][8] ) );
  FDN1QM1P \Queue_reg[0][8]  ( .D(n452), .CPN(Clk_r), .Q(Packet_Out[8]) );
  FDN1QM1P \Queue_reg[1][7]  ( .D(n419), .CPN(Clk_r), .Q(\Queue[1][7] ) );
  FDN1QM1P \Queue_reg[0][7]  ( .D(n451), .CPN(Clk_r), .Q(Packet_Out[7]) );
  FDN1QM1P \Queue_reg[1][6]  ( .D(n418), .CPN(Clk_r), .Q(\Queue[1][6] ) );
  FDN1QM1P \Queue_reg[0][6]  ( .D(n450), .CPN(Clk_r), .Q(Packet_Out[6]) );
  FDN1QM1P \Queue_reg[1][5]  ( .D(n417), .CPN(Clk_r), .Q(\Queue[1][5] ) );
  FDN1QM1P \Queue_reg[0][5]  ( .D(n449), .CPN(Clk_r), .Q(Packet_Out[5]) );
  FDN1QM1P \Queue_reg[1][4]  ( .D(n416), .CPN(Clk_r), .Q(\Queue[1][4] ) );
  FDN1QM1P \Queue_reg[0][4]  ( .D(n448), .CPN(Clk_r), .Q(Packet_Out[4]) );
  FDN1QM1P \Queue_reg[1][3]  ( .D(n415), .CPN(Clk_r), .Q(\Queue[1][3] ) );
  FDN1QM1P \Queue_reg[0][3]  ( .D(n447), .CPN(Clk_r), .Q(Packet_Out[3]) );
  FDN1QM1P \Queue_reg[1][2]  ( .D(n414), .CPN(Clk_r), .Q(\Queue[1][2] ) );
  FDN1QM1P \Queue_reg[0][2]  ( .D(n446), .CPN(Clk_r), .Q(Packet_Out[2]) );
  FDN1QM1P \Queue_reg[1][1]  ( .D(n413), .CPN(Clk_r), .Q(\Queue[1][1] ) );
  FDN1QM1P \Queue_reg[0][1]  ( .D(n445), .CPN(Clk_r), .Q(Packet_Out[1]) );
  FDN1QM1P \Queue_reg[1][0]  ( .D(n412), .CPN(Clk_r), .Q(\Queue[1][0] ) );
  FDN1QM1P \Queue_reg[0][0]  ( .D(n444), .CPN(Clk_r), .Q(Packet_Out[0]) );
  FDN2QM1P Empty_reg ( .D(n541), .CPN(Clk_r), .CD(Rst_n), .Q(n540) );
  BUFM2P U3 ( .A(n96), .Z(n6) );
  N1M2P U4 ( .A(n61), .Z(n93) );
  OAI211M4P U5 ( .A(n99), .B(n136), .C(Write_Ack), .D(n23), .Z(n58) );
  BUFM2P U6 ( .A(n131), .Z(n9) );
  BUFM2P U7 ( .A(n132), .Z(n10) );
  BUFM1P U8 ( .A(n131), .Z(n8) );
  AOI21M3P U9 ( .A(Write_Ack), .B(n141), .C(n140), .Z(n204) );
  NR3M1P U10 ( .A(Count[0]), .B(Count[2]), .C(n21), .Z(n99) );
  N1M1P U11 ( .A(n17), .Z(n138) );
  N1M1P U12 ( .A(Read_Ack), .Z(n136) );
  NR3M1P U13 ( .A(Count[2]), .B(n22), .C(n21), .Z(n139) );
  NR3M1P U14 ( .A(n22), .B(Count[2]), .C(Count[1]), .Z(n375) );
  OAI211M4P U15 ( .A(n139), .B(n136), .C(Write_Ack), .D(n97), .Z(n134) );
  OAI211M4P U16 ( .A(n141), .B(n136), .C(Write_Ack), .D(n135), .Z(n207) );
  OAI211M4P U17 ( .A(n139), .B(n138), .C(Rst_n), .D(n137), .Z(n205) );
  NR2FM3P U18 ( .A(n60), .B(n20), .Z(n19) );
  NR2M3P U19 ( .A(Read_Ack), .B(n98), .Z(n17) );
  NR3M1P U20 ( .A(Count[0]), .B(Count[1]), .C(n18), .Z(n141) );
  N1M3P U21 ( .A(Write_Ack), .Z(n98) );
  N1M1P U22 ( .A(n141), .Z(n20) );
  N1M1P U23 ( .A(Count[2]), .Z(n18) );
  N1M1P U24 ( .A(Count[1]), .Z(n21) );
  N1M1P U25 ( .A(Count[0]), .Z(n22) );
  OAI21M1P U26 ( .A(n60), .B(n59), .C(n140), .Z(n61) );
  ND2M2P U27 ( .A(n17), .B(Rst_n), .Z(n60) );
  AOI21M6P U28 ( .A(Write_Ack), .B(n99), .C(n140), .Z(n56) );
  ND2M2P U29 ( .A(Read_Ack), .B(Rst_n), .Z(n140) );
  AOI21M6P U30 ( .A(Write_Ack), .B(n375), .C(n140), .Z(n94) );
  N1M1P U31 ( .A(Packet_In[27]), .Z(n197) );
  N1M1P U32 ( .A(Packet_In[25]), .Z(n193) );
  N1M1P U33 ( .A(Packet_In[26]), .Z(n195) );
  N1M1P U34 ( .A(Packet_In[23]), .Z(n189) );
  N1M1P U35 ( .A(Packet_In[3]), .Z(n149) );
  N1M1P U36 ( .A(Packet_In[10]), .Z(n163) );
  N1M1P U37 ( .A(Packet_In[6]), .Z(n155) );
  N1M1P U38 ( .A(Packet_In[4]), .Z(n151) );
  N1M1P U39 ( .A(Packet_In[1]), .Z(n145) );
  N1M1P U40 ( .A(Packet_In[7]), .Z(n157) );
  N1M1P U41 ( .A(Packet_In[9]), .Z(n161) );
  N1M1P U42 ( .A(Packet_In[0]), .Z(n143) );
  N1M1P U43 ( .A(Packet_In[5]), .Z(n153) );
  N1M1P U44 ( .A(Packet_In[11]), .Z(n165) );
  N1M1P U45 ( .A(Packet_In[8]), .Z(n159) );
  N1M1P U46 ( .A(Packet_In[30]), .Z(n203) );
  N1M1P U47 ( .A(Packet_In[2]), .Z(n147) );
  N1M1P U48 ( .A(Packet_In[28]), .Z(n199) );
  N1M1P U49 ( .A(Packet_In[31]), .Z(n208) );
  N1M1P U50 ( .A(Packet_In[29]), .Z(n201) );
  N1M1P U51 ( .A(Packet_In[24]), .Z(n191) );
  N1M1P U52 ( .A(Packet_In[18]), .Z(n179) );
  N1M1P U53 ( .A(Packet_In[21]), .Z(n185) );
  N1M1P U54 ( .A(Packet_In[19]), .Z(n181) );
  N1M1P U55 ( .A(Packet_In[14]), .Z(n171) );
  N1M1P U56 ( .A(Packet_In[16]), .Z(n175) );
  N1M1P U57 ( .A(Packet_In[20]), .Z(n183) );
  N1M1P U58 ( .A(Packet_In[13]), .Z(n169) );
  N1M1P U59 ( .A(Packet_In[22]), .Z(n187) );
  N1M1P U60 ( .A(Packet_In[17]), .Z(n177) );
  N1M1P U61 ( .A(Packet_In[12]), .Z(n167) );
  N1M1P U62 ( .A(Packet_In[15]), .Z(n173) );
  BUFM2P U63 ( .A(n132), .Z(n11) );
  BUFM2P U64 ( .A(n55), .Z(n3) );
  BUFM2P U65 ( .A(n96), .Z(n7) );
  OAI211M1P U66 ( .A(n375), .B(n136), .C(Write_Ack), .D(n61), .Z(n96) );
  BUFM2P U67 ( .A(n55), .Z(n5) );
  BUFM2P U68 ( .A(n55), .Z(n4) );
  AOI22M1P U69 ( .A(Count[0]), .B(n138), .C(n16), .D(n22), .Z(n13) );
  OAI211M1P U70 ( .A(n99), .B(n138), .C(Rst_n), .D(n137), .Z(n132) );
  NR2M1P U71 ( .A(n136), .B(Write_Ack), .Z(n374) );
  NR2M1P U72 ( .A(n17), .B(n374), .Z(n373) );
  AOI22CDNM1P U73 ( .A(n373), .B(n22), .C(n373), .D(n22), .Z(n376) );
  N1M1P U74 ( .A(n374), .Z(n16) );
  AOI22CDNM1P U75 ( .A(Count[1]), .B(n13), .C(n13), .D(Count[1]), .Z(n377) );
  ND3M1P U76 ( .A(n22), .B(n18), .C(n21), .Z(n59) );
  ND2M1P U77 ( .A(Count[1]), .B(Read_Ack), .Z(n12) );
  OAI211M1P U78 ( .A(Count[1]), .B(n138), .C(n13), .D(n12), .Z(n14) );
  AOI22M1P U79 ( .A(n17), .B(n139), .C(Count[2]), .D(n14), .Z(n15) );
  OAI21M1P U80 ( .A(n59), .B(n16), .C(n15), .Z(n378) );
  AOI22CDNM1P U81 ( .A(n19), .B(n208), .C(\Queue[4][31] ), .D(n19), .Z(n379)
         );
  AOI22CDNM1P U82 ( .A(n19), .B(n143), .C(\Queue[4][0] ), .D(n19), .Z(n380) );
  AOI22CDNM1P U83 ( .A(n19), .B(n145), .C(\Queue[4][1] ), .D(n19), .Z(n381) );
  AOI22CDNM1P U84 ( .A(n19), .B(n147), .C(\Queue[4][2] ), .D(n19), .Z(n382) );
  AOI22CDNM1P U85 ( .A(n19), .B(n149), .C(\Queue[4][3] ), .D(n19), .Z(n383) );
  AOI22CDNM1P U86 ( .A(n19), .B(n151), .C(\Queue[4][4] ), .D(n19), .Z(n384) );
  AOI22CDNM1P U87 ( .A(n19), .B(n153), .C(\Queue[4][5] ), .D(n19), .Z(n385) );
  AOI22CDNM1P U88 ( .A(n19), .B(n155), .C(\Queue[4][6] ), .D(n19), .Z(n386) );
  AOI22CDNM1P U89 ( .A(n19), .B(n157), .C(\Queue[4][7] ), .D(n19), .Z(n387) );
  AOI22CDNM1P U90 ( .A(n19), .B(n159), .C(\Queue[4][8] ), .D(n19), .Z(n388) );
  AOI22CDNM1P U91 ( .A(n19), .B(n161), .C(\Queue[4][9] ), .D(n19), .Z(n389) );
  AOI22CDNM1P U92 ( .A(n19), .B(n163), .C(\Queue[4][10] ), .D(n19), .Z(n390)
         );
  AOI22CDNM1P U93 ( .A(n19), .B(n165), .C(\Queue[4][11] ), .D(n19), .Z(n391)
         );
  AOI22CDNM1P U94 ( .A(n19), .B(n167), .C(\Queue[4][12] ), .D(n19), .Z(n392)
         );
  AOI22CDNM1P U95 ( .A(n19), .B(n169), .C(\Queue[4][13] ), .D(n19), .Z(n393)
         );
  AOI22CDNM1P U96 ( .A(n19), .B(n171), .C(\Queue[4][14] ), .D(n19), .Z(n394)
         );
  AOI22CDNM1P U97 ( .A(n19), .B(n173), .C(\Queue[4][15] ), .D(n19), .Z(n395)
         );
  AOI22CDNM1P U98 ( .A(n19), .B(n175), .C(\Queue[4][16] ), .D(n19), .Z(n396)
         );
  AOI22CDNM1P U99 ( .A(n19), .B(n177), .C(\Queue[4][17] ), .D(n19), .Z(n397)
         );
  AOI22CDNM1P U100 ( .A(n19), .B(n179), .C(\Queue[4][18] ), .D(n19), .Z(n398)
         );
  AOI22CDNM1P U101 ( .A(n19), .B(n181), .C(\Queue[4][19] ), .D(n19), .Z(n399)
         );
  AOI22CDNM1P U102 ( .A(n19), .B(n183), .C(\Queue[4][20] ), .D(n19), .Z(n400)
         );
  AOI22CDNM1P U103 ( .A(n19), .B(n185), .C(\Queue[4][21] ), .D(n19), .Z(n401)
         );
  AOI22CDNM1P U104 ( .A(n19), .B(n187), .C(\Queue[4][22] ), .D(n19), .Z(n402)
         );
  AOI22CDNM1P U105 ( .A(n19), .B(n189), .C(\Queue[4][23] ), .D(n19), .Z(n403)
         );
  AOI22CDNM1P U106 ( .A(n19), .B(n191), .C(\Queue[4][24] ), .D(n19), .Z(n404)
         );
  AOI22CDNM1P U107 ( .A(n19), .B(n193), .C(\Queue[4][25] ), .D(n19), .Z(n405)
         );
  AOI22CDNM1P U108 ( .A(n19), .B(n195), .C(\Queue[4][26] ), .D(n19), .Z(n406)
         );
  AOI22CDNM1P U109 ( .A(n19), .B(n197), .C(\Queue[4][27] ), .D(n19), .Z(n407)
         );
  AOI22CDNM1P U110 ( .A(n19), .B(n199), .C(\Queue[4][28] ), .D(n19), .Z(n408)
         );
  AOI22CDNM1P U111 ( .A(n19), .B(n201), .C(\Queue[4][29] ), .D(n19), .Z(n409)
         );
  AOI22CDNM1P U112 ( .A(n19), .B(n203), .C(\Queue[4][30] ), .D(n19), .Z(n410)
         );
  OAI22CDNM1P U113 ( .A(n138), .B(n20), .C(n373), .D(Full), .Z(n411) );
  OA21M1P U114 ( .A(n138), .B(n375), .C(Rst_n), .Z(n23) );
  OAI21M1P U115 ( .A(Write_Ack), .B(Read_Ack), .C(n23), .Z(n55) );
  AOI22M1P U116 ( .A(\Queue[2][0] ), .B(n56), .C(\Queue[1][0] ), .D(n3), .Z(
        n24) );
  OAI21M1P U117 ( .A(n143), .B(n58), .C(n24), .Z(n412) );
  AOI22M1P U118 ( .A(n56), .B(\Queue[2][1] ), .C(\Queue[1][1] ), .D(n3), .Z(
        n25) );
  OAI21M1P U119 ( .A(n58), .B(n145), .C(n25), .Z(n413) );
  AOI22M1P U120 ( .A(n56), .B(\Queue[2][2] ), .C(\Queue[1][2] ), .D(n3), .Z(
        n26) );
  OAI21M1P U121 ( .A(n58), .B(n147), .C(n26), .Z(n414) );
  AOI22M1P U122 ( .A(n56), .B(\Queue[2][3] ), .C(\Queue[1][3] ), .D(n3), .Z(
        n27) );
  OAI21M1P U123 ( .A(n58), .B(n149), .C(n27), .Z(n415) );
  AOI22M1P U124 ( .A(n56), .B(\Queue[2][4] ), .C(\Queue[1][4] ), .D(n3), .Z(
        n28) );
  OAI21M1P U125 ( .A(n58), .B(n151), .C(n28), .Z(n416) );
  AOI22M1P U126 ( .A(n56), .B(\Queue[2][5] ), .C(\Queue[1][5] ), .D(n3), .Z(
        n29) );
  OAI21M1P U127 ( .A(n58), .B(n153), .C(n29), .Z(n417) );
  AOI22M1P U128 ( .A(n56), .B(\Queue[2][6] ), .C(\Queue[1][6] ), .D(n3), .Z(
        n30) );
  OAI21M1P U129 ( .A(n58), .B(n155), .C(n30), .Z(n418) );
  AOI22M1P U130 ( .A(n56), .B(\Queue[2][7] ), .C(\Queue[1][7] ), .D(n3), .Z(
        n31) );
  OAI21M1P U131 ( .A(n58), .B(n157), .C(n31), .Z(n419) );
  AOI22M1P U132 ( .A(n56), .B(\Queue[2][8] ), .C(\Queue[1][8] ), .D(n3), .Z(
        n32) );
  OAI21M1P U133 ( .A(n58), .B(n159), .C(n32), .Z(n420) );
  AOI22M1P U134 ( .A(n56), .B(\Queue[2][9] ), .C(\Queue[1][9] ), .D(n4), .Z(
        n33) );
  OAI21M1P U135 ( .A(n58), .B(n161), .C(n33), .Z(n421) );
  AOI22M1P U136 ( .A(n56), .B(\Queue[2][10] ), .C(\Queue[1][10] ), .D(n4), .Z(
        n34) );
  OAI21M1P U137 ( .A(n58), .B(n163), .C(n34), .Z(n422) );
  AOI22M1P U138 ( .A(n56), .B(\Queue[2][11] ), .C(\Queue[1][11] ), .D(n4), .Z(
        n35) );
  OAI21M1P U139 ( .A(n58), .B(n165), .C(n35), .Z(n423) );
  AOI22M1P U140 ( .A(n56), .B(\Queue[2][12] ), .C(\Queue[1][12] ), .D(n4), .Z(
        n36) );
  OAI21M1P U141 ( .A(n58), .B(n167), .C(n36), .Z(n424) );
  AOI22M1P U142 ( .A(n56), .B(\Queue[2][13] ), .C(\Queue[1][13] ), .D(n4), .Z(
        n37) );
  OAI21M1P U143 ( .A(n58), .B(n169), .C(n37), .Z(n425) );
  AOI22M1P U144 ( .A(n56), .B(\Queue[2][14] ), .C(\Queue[1][14] ), .D(n4), .Z(
        n38) );
  OAI21M1P U145 ( .A(n58), .B(n171), .C(n38), .Z(n426) );
  AOI22M1P U146 ( .A(n56), .B(\Queue[2][15] ), .C(\Queue[1][15] ), .D(n4), .Z(
        n39) );
  OAI21M1P U147 ( .A(n58), .B(n173), .C(n39), .Z(n427) );
  AOI22M1P U148 ( .A(n56), .B(\Queue[2][16] ), .C(\Queue[1][16] ), .D(n4), .Z(
        n40) );
  OAI21M1P U149 ( .A(n58), .B(n175), .C(n40), .Z(n428) );
  AOI22M1P U150 ( .A(n56), .B(\Queue[2][17] ), .C(\Queue[1][17] ), .D(n4), .Z(
        n41) );
  OAI21M1P U151 ( .A(n58), .B(n177), .C(n41), .Z(n429) );
  AOI22M1P U152 ( .A(n56), .B(\Queue[2][18] ), .C(\Queue[1][18] ), .D(n5), .Z(
        n42) );
  OAI21M1P U153 ( .A(n58), .B(n179), .C(n42), .Z(n430) );
  AOI22M1P U154 ( .A(n56), .B(\Queue[2][19] ), .C(\Queue[1][19] ), .D(n5), .Z(
        n43) );
  OAI21M1P U155 ( .A(n58), .B(n181), .C(n43), .Z(n431) );
  AOI22M1P U156 ( .A(n56), .B(\Queue[2][20] ), .C(\Queue[1][20] ), .D(n5), .Z(
        n44) );
  OAI21M1P U157 ( .A(n58), .B(n183), .C(n44), .Z(n432) );
  AOI22M1P U158 ( .A(n56), .B(\Queue[2][21] ), .C(\Queue[1][21] ), .D(n5), .Z(
        n45) );
  OAI21M1P U159 ( .A(n58), .B(n185), .C(n45), .Z(n433) );
  AOI22M1P U160 ( .A(n56), .B(\Queue[2][22] ), .C(\Queue[1][22] ), .D(n5), .Z(
        n46) );
  OAI21M1P U161 ( .A(n58), .B(n187), .C(n46), .Z(n434) );
  AOI22M1P U162 ( .A(n56), .B(\Queue[2][23] ), .C(\Queue[1][23] ), .D(n5), .Z(
        n47) );
  OAI21M1P U163 ( .A(n58), .B(n189), .C(n47), .Z(n435) );
  AOI22M1P U164 ( .A(n56), .B(\Queue[2][24] ), .C(\Queue[1][24] ), .D(n5), .Z(
        n48) );
  OAI21M1P U165 ( .A(n58), .B(n191), .C(n48), .Z(n436) );
  AOI22M1P U166 ( .A(n56), .B(\Queue[2][25] ), .C(\Queue[1][25] ), .D(n5), .Z(
        n49) );
  OAI21M1P U167 ( .A(n58), .B(n193), .C(n49), .Z(n437) );
  AOI22M1P U168 ( .A(n56), .B(\Queue[2][26] ), .C(\Queue[1][26] ), .D(n5), .Z(
        n50) );
  OAI21M1P U169 ( .A(n58), .B(n195), .C(n50), .Z(n438) );
  AOI22M1P U170 ( .A(n56), .B(\Queue[2][27] ), .C(\Queue[1][27] ), .D(n3), .Z(
        n51) );
  OAI21M1P U171 ( .A(n58), .B(n197), .C(n51), .Z(n439) );
  AOI22M1P U172 ( .A(n56), .B(\Queue[2][28] ), .C(\Queue[1][28] ), .D(n4), .Z(
        n52) );
  OAI21M1P U173 ( .A(n58), .B(n199), .C(n52), .Z(n440) );
  AOI22M1P U174 ( .A(n56), .B(\Queue[2][29] ), .C(\Queue[1][29] ), .D(n5), .Z(
        n53) );
  OAI21M1P U175 ( .A(n58), .B(n201), .C(n53), .Z(n441) );
  AOI22M1P U176 ( .A(n56), .B(\Queue[2][30] ), .C(\Queue[1][30] ), .D(n4), .Z(
        n54) );
  OAI21M1P U177 ( .A(n58), .B(n203), .C(n54), .Z(n442) );
  AOI22M1P U178 ( .A(n56), .B(\Queue[2][31] ), .C(\Queue[1][31] ), .D(n5), .Z(
        n57) );
  OAI21M1P U179 ( .A(n58), .B(n208), .C(n57), .Z(n443) );
  AOI22M1P U180 ( .A(\Queue[1][0] ), .B(n94), .C(n93), .D(Packet_Out[0]), .Z(
        n62) );
  OAI21M1P U181 ( .A(n143), .B(n6), .C(n62), .Z(n444) );
  AOI22M1P U182 ( .A(\Queue[1][1] ), .B(n94), .C(n93), .D(Packet_Out[1]), .Z(
        n63) );
  OAI21M1P U183 ( .A(n145), .B(n6), .C(n63), .Z(n445) );
  AOI22M1P U184 ( .A(\Queue[1][2] ), .B(n94), .C(n93), .D(Packet_Out[2]), .Z(
        n64) );
  OAI21M1P U185 ( .A(n147), .B(n6), .C(n64), .Z(n446) );
  AOI22M1P U186 ( .A(\Queue[1][3] ), .B(n94), .C(n93), .D(Packet_Out[3]), .Z(
        n65) );
  OAI21M1P U187 ( .A(n149), .B(n6), .C(n65), .Z(n447) );
  AOI22M1P U188 ( .A(\Queue[1][4] ), .B(n94), .C(n93), .D(Packet_Out[4]), .Z(
        n66) );
  OAI21M1P U189 ( .A(n151), .B(n6), .C(n66), .Z(n448) );
  AOI22M1P U190 ( .A(\Queue[1][5] ), .B(n94), .C(n93), .D(Packet_Out[5]), .Z(
        n67) );
  OAI21M1P U191 ( .A(n153), .B(n6), .C(n67), .Z(n449) );
  AOI22M1P U192 ( .A(\Queue[1][6] ), .B(n94), .C(n93), .D(Packet_Out[6]), .Z(
        n68) );
  OAI21M1P U193 ( .A(n155), .B(n6), .C(n68), .Z(n450) );
  AOI22M1P U194 ( .A(\Queue[1][7] ), .B(n94), .C(n93), .D(Packet_Out[7]), .Z(
        n69) );
  OAI21M1P U195 ( .A(n157), .B(n6), .C(n69), .Z(n451) );
  AOI22M1P U196 ( .A(\Queue[1][8] ), .B(n94), .C(n93), .D(Packet_Out[8]), .Z(
        n70) );
  OAI21M1P U197 ( .A(n159), .B(n6), .C(n70), .Z(n452) );
  AOI22M1P U198 ( .A(\Queue[1][9] ), .B(n94), .C(n93), .D(Packet_Out[9]), .Z(
        n71) );
  OAI21M1P U199 ( .A(n161), .B(n6), .C(n71), .Z(n453) );
  AOI22M1P U200 ( .A(\Queue[1][10] ), .B(n94), .C(n93), .D(Packet_Out[10]), 
        .Z(n72) );
  OAI21M1P U201 ( .A(n163), .B(n6), .C(n72), .Z(n454) );
  AOI22M1P U202 ( .A(\Queue[1][11] ), .B(n94), .C(n93), .D(Packet_Out[11]), 
        .Z(n73) );
  OAI21M1P U203 ( .A(n165), .B(n6), .C(n73), .Z(n455) );
  AOI22M1P U204 ( .A(\Queue[1][12] ), .B(n94), .C(n93), .D(Packet_Out[12]), 
        .Z(n74) );
  OAI21M1P U205 ( .A(n167), .B(n6), .C(n74), .Z(n456) );
  AOI22M1P U206 ( .A(\Queue[1][13] ), .B(n94), .C(n93), .D(Packet_Out[13]), 
        .Z(n75) );
  OAI21M1P U207 ( .A(n169), .B(n6), .C(n75), .Z(n457) );
  AOI22M1P U208 ( .A(\Queue[1][14] ), .B(n94), .C(n93), .D(Packet_Out[14]), 
        .Z(n76) );
  OAI21M1P U209 ( .A(n171), .B(n6), .C(n76), .Z(n458) );
  AOI22M1P U210 ( .A(\Queue[1][15] ), .B(n94), .C(n93), .D(Packet_Out[15]), 
        .Z(n77) );
  OAI21M1P U211 ( .A(n173), .B(n6), .C(n77), .Z(n459) );
  AOI22M1P U212 ( .A(\Queue[1][16] ), .B(n94), .C(n93), .D(Packet_Out[16]), 
        .Z(n78) );
  OAI21M1P U213 ( .A(n175), .B(n6), .C(n78), .Z(n460) );
  AOI22M1P U214 ( .A(\Queue[1][17] ), .B(n94), .C(n93), .D(Packet_Out[17]), 
        .Z(n79) );
  OAI21M1P U215 ( .A(n177), .B(n6), .C(n79), .Z(n461) );
  AOI22M1P U216 ( .A(\Queue[1][18] ), .B(n94), .C(n93), .D(Packet_Out[18]), 
        .Z(n80) );
  OAI21M1P U217 ( .A(n179), .B(n6), .C(n80), .Z(n462) );
  AOI22M1P U218 ( .A(\Queue[1][19] ), .B(n94), .C(n93), .D(Packet_Out[19]), 
        .Z(n81) );
  OAI21M1P U219 ( .A(n181), .B(n6), .C(n81), .Z(n463) );
  AOI22M1P U220 ( .A(\Queue[1][20] ), .B(n94), .C(n93), .D(Packet_Out[20]), 
        .Z(n82) );
  OAI21M1P U221 ( .A(n183), .B(n7), .C(n82), .Z(n464) );
  AOI22M1P U222 ( .A(\Queue[1][21] ), .B(n94), .C(n93), .D(Packet_Out[21]), 
        .Z(n83) );
  OAI21M1P U223 ( .A(n185), .B(n7), .C(n83), .Z(n465) );
  AOI22M1P U224 ( .A(\Queue[1][22] ), .B(n94), .C(n93), .D(Packet_Out[22]), 
        .Z(n84) );
  OAI21M1P U225 ( .A(n187), .B(n7), .C(n84), .Z(n466) );
  AOI22M1P U226 ( .A(\Queue[1][23] ), .B(n94), .C(n93), .D(Packet_Out[23]), 
        .Z(n85) );
  OAI21M1P U227 ( .A(n189), .B(n7), .C(n85), .Z(n467) );
  AOI22M1P U228 ( .A(\Queue[1][24] ), .B(n94), .C(n93), .D(Packet_Out[24]), 
        .Z(n86) );
  OAI21M1P U229 ( .A(n191), .B(n7), .C(n86), .Z(n468) );
  AOI22M1P U230 ( .A(\Queue[1][25] ), .B(n94), .C(n93), .D(Packet_Out[25]), 
        .Z(n87) );
  OAI21M1P U231 ( .A(n193), .B(n7), .C(n87), .Z(n469) );
  AOI22M1P U232 ( .A(\Queue[1][26] ), .B(n94), .C(n93), .D(Packet_Out[26]), 
        .Z(n88) );
  OAI21M1P U233 ( .A(n195), .B(n7), .C(n88), .Z(n470) );
  AOI22M1P U234 ( .A(\Queue[1][27] ), .B(n94), .C(n93), .D(Packet_Out[27]), 
        .Z(n89) );
  OAI21M1P U235 ( .A(n197), .B(n7), .C(n89), .Z(n471) );
  AOI22M1P U236 ( .A(\Queue[1][28] ), .B(n94), .C(n93), .D(Packet_Out[28]), 
        .Z(n90) );
  OAI21M1P U237 ( .A(n199), .B(n7), .C(n90), .Z(n472) );
  AOI22M1P U238 ( .A(\Queue[1][29] ), .B(n94), .C(n93), .D(Packet_Out[29]), 
        .Z(n91) );
  OAI21M1P U239 ( .A(n201), .B(n7), .C(n91), .Z(n473) );
  AOI22M1P U240 ( .A(\Queue[1][30] ), .B(n94), .C(n93), .D(Packet_Out[30]), 
        .Z(n92) );
  OAI21M1P U241 ( .A(n203), .B(n6), .C(n92), .Z(n474) );
  AOI22M1P U242 ( .A(\Queue[1][31] ), .B(n94), .C(n93), .D(Packet_Out[31]), 
        .Z(n95) );
  OAI21M1P U243 ( .A(n208), .B(n7), .C(n95), .Z(n475) );
  OA21M1P U244 ( .A(n138), .B(n99), .C(Rst_n), .Z(n97) );
  ND2M1P U245 ( .A(n98), .B(n136), .Z(n137) );
  AOI21M1P U246 ( .A(Write_Ack), .B(n139), .C(n140), .Z(n131) );
  AOI22M1P U247 ( .A(\Queue[2][0] ), .B(n10), .C(\Queue[3][0] ), .D(n8), .Z(
        n100) );
  OAI21M1P U248 ( .A(n143), .B(n134), .C(n100), .Z(n476) );
  AOI22M1P U249 ( .A(\Queue[2][1] ), .B(n10), .C(n9), .D(\Queue[3][1] ), .Z(
        n101) );
  OAI21M1P U250 ( .A(n145), .B(n134), .C(n101), .Z(n477) );
  AOI22M1P U251 ( .A(\Queue[2][2] ), .B(n10), .C(n9), .D(\Queue[3][2] ), .Z(
        n102) );
  OAI21M1P U252 ( .A(n147), .B(n134), .C(n102), .Z(n478) );
  AOI22M1P U253 ( .A(\Queue[2][3] ), .B(n10), .C(n9), .D(\Queue[3][3] ), .Z(
        n103) );
  OAI21M1P U254 ( .A(n149), .B(n134), .C(n103), .Z(n479) );
  AOI22M1P U255 ( .A(\Queue[2][4] ), .B(n10), .C(n9), .D(\Queue[3][4] ), .Z(
        n104) );
  OAI21M1P U256 ( .A(n151), .B(n134), .C(n104), .Z(n480) );
  AOI22M1P U257 ( .A(\Queue[2][5] ), .B(n10), .C(n9), .D(\Queue[3][5] ), .Z(
        n105) );
  OAI21M1P U258 ( .A(n153), .B(n134), .C(n105), .Z(n481) );
  AOI22M1P U259 ( .A(\Queue[2][6] ), .B(n10), .C(n9), .D(\Queue[3][6] ), .Z(
        n106) );
  OAI21M1P U260 ( .A(n155), .B(n134), .C(n106), .Z(n482) );
  AOI22M1P U261 ( .A(\Queue[2][7] ), .B(n10), .C(n9), .D(\Queue[3][7] ), .Z(
        n107) );
  OAI21M1P U262 ( .A(n157), .B(n134), .C(n107), .Z(n483) );
  AOI22M1P U263 ( .A(\Queue[2][8] ), .B(n10), .C(n9), .D(\Queue[3][8] ), .Z(
        n108) );
  OAI21M1P U264 ( .A(n159), .B(n134), .C(n108), .Z(n484) );
  AOI22M1P U265 ( .A(\Queue[2][9] ), .B(n10), .C(n9), .D(\Queue[3][9] ), .Z(
        n109) );
  OAI21M1P U266 ( .A(n161), .B(n134), .C(n109), .Z(n485) );
  AOI22M1P U267 ( .A(\Queue[2][10] ), .B(n10), .C(n9), .D(\Queue[3][10] ), .Z(
        n110) );
  OAI21M1P U268 ( .A(n163), .B(n134), .C(n110), .Z(n486) );
  AOI22M1P U269 ( .A(\Queue[2][11] ), .B(n10), .C(n9), .D(\Queue[3][11] ), .Z(
        n111) );
  OAI21M1P U270 ( .A(n165), .B(n134), .C(n111), .Z(n487) );
  AOI22M1P U271 ( .A(\Queue[2][12] ), .B(n10), .C(n9), .D(\Queue[3][12] ), .Z(
        n112) );
  OAI21M1P U272 ( .A(n167), .B(n134), .C(n112), .Z(n488) );
  AOI22M1P U273 ( .A(\Queue[2][13] ), .B(n10), .C(n9), .D(\Queue[3][13] ), .Z(
        n113) );
  OAI21M1P U274 ( .A(n169), .B(n134), .C(n113), .Z(n489) );
  AOI22M1P U275 ( .A(\Queue[2][14] ), .B(n10), .C(n9), .D(\Queue[3][14] ), .Z(
        n114) );
  OAI21M1P U276 ( .A(n171), .B(n134), .C(n114), .Z(n490) );
  AOI22M1P U277 ( .A(\Queue[2][15] ), .B(n10), .C(n9), .D(\Queue[3][15] ), .Z(
        n115) );
  OAI21M1P U278 ( .A(n173), .B(n134), .C(n115), .Z(n491) );
  AOI22M1P U279 ( .A(\Queue[2][16] ), .B(n10), .C(n9), .D(\Queue[3][16] ), .Z(
        n116) );
  OAI21M1P U280 ( .A(n175), .B(n134), .C(n116), .Z(n492) );
  AOI22M1P U281 ( .A(\Queue[2][17] ), .B(n10), .C(n9), .D(\Queue[3][17] ), .Z(
        n117) );
  OAI21M1P U282 ( .A(n177), .B(n134), .C(n117), .Z(n493) );
  AOI22M1P U283 ( .A(\Queue[2][18] ), .B(n10), .C(n9), .D(\Queue[3][18] ), .Z(
        n118) );
  OAI21M1P U284 ( .A(n179), .B(n134), .C(n118), .Z(n494) );
  AOI22M1P U285 ( .A(\Queue[2][19] ), .B(n10), .C(n9), .D(\Queue[3][19] ), .Z(
        n119) );
  OAI21M1P U286 ( .A(n181), .B(n134), .C(n119), .Z(n495) );
  AOI22M1P U287 ( .A(\Queue[2][20] ), .B(n11), .C(n9), .D(\Queue[3][20] ), .Z(
        n120) );
  OAI21M1P U288 ( .A(n183), .B(n134), .C(n120), .Z(n496) );
  AOI22M1P U289 ( .A(\Queue[2][21] ), .B(n11), .C(n9), .D(\Queue[3][21] ), .Z(
        n121) );
  OAI21M1P U290 ( .A(n185), .B(n134), .C(n121), .Z(n497) );
  AOI22M1P U291 ( .A(\Queue[2][22] ), .B(n11), .C(n8), .D(\Queue[3][22] ), .Z(
        n122) );
  OAI21M1P U292 ( .A(n187), .B(n134), .C(n122), .Z(n498) );
  AOI22M1P U293 ( .A(\Queue[2][23] ), .B(n11), .C(n8), .D(\Queue[3][23] ), .Z(
        n123) );
  OAI21M1P U294 ( .A(n189), .B(n134), .C(n123), .Z(n499) );
  AOI22M1P U295 ( .A(\Queue[2][24] ), .B(n11), .C(n8), .D(\Queue[3][24] ), .Z(
        n124) );
  OAI21M1P U296 ( .A(n191), .B(n134), .C(n124), .Z(n500) );
  AOI22M1P U297 ( .A(\Queue[2][25] ), .B(n11), .C(n8), .D(\Queue[3][25] ), .Z(
        n125) );
  OAI21M1P U298 ( .A(n193), .B(n134), .C(n125), .Z(n501) );
  AOI22M1P U299 ( .A(\Queue[2][26] ), .B(n11), .C(n8), .D(\Queue[3][26] ), .Z(
        n126) );
  OAI21M1P U300 ( .A(n195), .B(n134), .C(n126), .Z(n502) );
  AOI22M1P U301 ( .A(\Queue[2][27] ), .B(n11), .C(n8), .D(\Queue[3][27] ), .Z(
        n127) );
  OAI21M1P U302 ( .A(n197), .B(n134), .C(n127), .Z(n503) );
  AOI22M1P U303 ( .A(\Queue[2][28] ), .B(n11), .C(n8), .D(\Queue[3][28] ), .Z(
        n128) );
  OAI21M1P U304 ( .A(n199), .B(n134), .C(n128), .Z(n504) );
  AOI22M1P U305 ( .A(\Queue[2][29] ), .B(n11), .C(n8), .D(\Queue[3][29] ), .Z(
        n129) );
  OAI21M1P U306 ( .A(n201), .B(n134), .C(n129), .Z(n505) );
  AOI22M1P U307 ( .A(\Queue[2][30] ), .B(n10), .C(n8), .D(\Queue[3][30] ), .Z(
        n130) );
  OAI21M1P U308 ( .A(n203), .B(n134), .C(n130), .Z(n506) );
  AOI22M1P U309 ( .A(\Queue[2][31] ), .B(n11), .C(n8), .D(\Queue[3][31] ), .Z(
        n133) );
  OAI21M1P U310 ( .A(n208), .B(n134), .C(n133), .Z(n507) );
  OA21M1P U311 ( .A(n138), .B(n139), .C(Rst_n), .Z(n135) );
  AOI22M1P U312 ( .A(\Queue[3][0] ), .B(n205), .C(n204), .D(\Queue[4][0] ), 
        .Z(n142) );
  OAI21M1P U313 ( .A(n143), .B(n207), .C(n142), .Z(n508) );
  AOI22M1P U314 ( .A(\Queue[3][1] ), .B(n205), .C(n204), .D(\Queue[4][1] ), 
        .Z(n144) );
  OAI21M1P U315 ( .A(n145), .B(n207), .C(n144), .Z(n509) );
  AOI22M1P U316 ( .A(\Queue[3][2] ), .B(n205), .C(n204), .D(\Queue[4][2] ), 
        .Z(n146) );
  OAI21M1P U317 ( .A(n147), .B(n207), .C(n146), .Z(n510) );
  AOI22M1P U318 ( .A(\Queue[3][3] ), .B(n205), .C(n204), .D(\Queue[4][3] ), 
        .Z(n148) );
  OAI21M1P U319 ( .A(n149), .B(n207), .C(n148), .Z(n511) );
  AOI22M1P U320 ( .A(\Queue[3][4] ), .B(n205), .C(n204), .D(\Queue[4][4] ), 
        .Z(n150) );
  OAI21M1P U321 ( .A(n151), .B(n207), .C(n150), .Z(n512) );
  AOI22M1P U322 ( .A(\Queue[3][5] ), .B(n205), .C(n204), .D(\Queue[4][5] ), 
        .Z(n152) );
  OAI21M1P U323 ( .A(n153), .B(n207), .C(n152), .Z(n513) );
  AOI22M1P U324 ( .A(\Queue[3][6] ), .B(n205), .C(n204), .D(\Queue[4][6] ), 
        .Z(n154) );
  OAI21M1P U325 ( .A(n155), .B(n207), .C(n154), .Z(n514) );
  AOI22M1P U326 ( .A(\Queue[3][7] ), .B(n205), .C(n204), .D(\Queue[4][7] ), 
        .Z(n156) );
  OAI21M1P U327 ( .A(n157), .B(n207), .C(n156), .Z(n515) );
  AOI22M1P U328 ( .A(\Queue[3][8] ), .B(n205), .C(n204), .D(\Queue[4][8] ), 
        .Z(n158) );
  OAI21M1P U329 ( .A(n159), .B(n207), .C(n158), .Z(n516) );
  AOI22M1P U330 ( .A(\Queue[3][9] ), .B(n205), .C(n204), .D(\Queue[4][9] ), 
        .Z(n160) );
  OAI21M1P U331 ( .A(n161), .B(n207), .C(n160), .Z(n517) );
  AOI22M1P U332 ( .A(\Queue[3][10] ), .B(n205), .C(n204), .D(\Queue[4][10] ), 
        .Z(n162) );
  OAI21M1P U333 ( .A(n163), .B(n207), .C(n162), .Z(n518) );
  AOI22M1P U334 ( .A(\Queue[3][11] ), .B(n205), .C(n204), .D(\Queue[4][11] ), 
        .Z(n164) );
  OAI21M1P U335 ( .A(n165), .B(n207), .C(n164), .Z(n519) );
  AOI22M1P U336 ( .A(\Queue[3][12] ), .B(n205), .C(n204), .D(\Queue[4][12] ), 
        .Z(n166) );
  OAI21M1P U337 ( .A(n167), .B(n207), .C(n166), .Z(n520) );
  AOI22M1P U338 ( .A(\Queue[3][13] ), .B(n205), .C(n204), .D(\Queue[4][13] ), 
        .Z(n168) );
  OAI21M1P U339 ( .A(n169), .B(n207), .C(n168), .Z(n521) );
  AOI22M1P U340 ( .A(\Queue[3][14] ), .B(n205), .C(n204), .D(\Queue[4][14] ), 
        .Z(n170) );
  OAI21M1P U341 ( .A(n171), .B(n207), .C(n170), .Z(n522) );
  AOI22M1P U342 ( .A(\Queue[3][15] ), .B(n205), .C(n204), .D(\Queue[4][15] ), 
        .Z(n172) );
  OAI21M1P U343 ( .A(n173), .B(n207), .C(n172), .Z(n523) );
  AOI22M1P U344 ( .A(\Queue[3][16] ), .B(n205), .C(n204), .D(\Queue[4][16] ), 
        .Z(n174) );
  OAI21M1P U345 ( .A(n175), .B(n207), .C(n174), .Z(n524) );
  AOI22M1P U346 ( .A(\Queue[3][17] ), .B(n205), .C(n204), .D(\Queue[4][17] ), 
        .Z(n176) );
  OAI21M1P U347 ( .A(n177), .B(n207), .C(n176), .Z(n525) );
  AOI22M1P U348 ( .A(\Queue[3][18] ), .B(n205), .C(n204), .D(\Queue[4][18] ), 
        .Z(n178) );
  OAI21M1P U349 ( .A(n179), .B(n207), .C(n178), .Z(n526) );
  AOI22M1P U350 ( .A(\Queue[3][19] ), .B(n205), .C(n204), .D(\Queue[4][19] ), 
        .Z(n180) );
  OAI21M1P U351 ( .A(n181), .B(n207), .C(n180), .Z(n527) );
  AOI22M1P U352 ( .A(\Queue[3][20] ), .B(n205), .C(n204), .D(\Queue[4][20] ), 
        .Z(n182) );
  OAI21M1P U353 ( .A(n183), .B(n207), .C(n182), .Z(n528) );
  AOI22M1P U354 ( .A(\Queue[3][21] ), .B(n205), .C(n204), .D(\Queue[4][21] ), 
        .Z(n184) );
  OAI21M1P U355 ( .A(n185), .B(n207), .C(n184), .Z(n529) );
  AOI22M1P U356 ( .A(\Queue[3][22] ), .B(n205), .C(n204), .D(\Queue[4][22] ), 
        .Z(n186) );
  OAI21M1P U357 ( .A(n187), .B(n207), .C(n186), .Z(n530) );
  AOI22M1P U358 ( .A(\Queue[3][23] ), .B(n205), .C(n204), .D(\Queue[4][23] ), 
        .Z(n188) );
  OAI21M1P U359 ( .A(n189), .B(n207), .C(n188), .Z(n531) );
  AOI22M1P U360 ( .A(\Queue[3][24] ), .B(n205), .C(n204), .D(\Queue[4][24] ), 
        .Z(n190) );
  OAI21M1P U361 ( .A(n191), .B(n207), .C(n190), .Z(n532) );
  AOI22M1P U362 ( .A(\Queue[3][25] ), .B(n205), .C(n204), .D(\Queue[4][25] ), 
        .Z(n192) );
  OAI21M1P U363 ( .A(n193), .B(n207), .C(n192), .Z(n533) );
  AOI22M1P U364 ( .A(\Queue[3][26] ), .B(n205), .C(n204), .D(\Queue[4][26] ), 
        .Z(n194) );
  OAI21M1P U365 ( .A(n195), .B(n207), .C(n194), .Z(n534) );
  AOI22M1P U366 ( .A(\Queue[3][27] ), .B(n205), .C(n204), .D(\Queue[4][27] ), 
        .Z(n196) );
  OAI21M1P U367 ( .A(n197), .B(n207), .C(n196), .Z(n535) );
  AOI22M1P U368 ( .A(\Queue[3][28] ), .B(n205), .C(n204), .D(\Queue[4][28] ), 
        .Z(n198) );
  OAI21M1P U369 ( .A(n199), .B(n207), .C(n198), .Z(n536) );
  AOI22M1P U370 ( .A(\Queue[3][29] ), .B(n205), .C(n204), .D(\Queue[4][29] ), 
        .Z(n200) );
  OAI21M1P U371 ( .A(n201), .B(n207), .C(n200), .Z(n537) );
  AOI22M1P U372 ( .A(\Queue[3][30] ), .B(n205), .C(n204), .D(\Queue[4][30] ), 
        .Z(n202) );
  OAI21M1P U373 ( .A(n203), .B(n207), .C(n202), .Z(n538) );
  AOI22M1P U374 ( .A(\Queue[3][31] ), .B(n205), .C(n204), .D(\Queue[4][31] ), 
        .Z(n206) );
  OAI21M1P U375 ( .A(n208), .B(n207), .C(n206), .Z(n539) );
  N1M1P U376 ( .A(n540), .Z(Empty) );
  AOI22M1P U377 ( .A(n375), .B(n374), .C(n373), .D(Empty), .Z(n541) );
endmodule


module Packet_Queue_6 ( Clk_r, Rst_n, Packet_In, Read_Ack, Write_Ack, 
        Packet_Out, Empty, Full );
  input [31:0] Packet_In;
  output [31:0] Packet_Out;
  input Clk_r, Rst_n, Read_Ack, Write_Ack;
  output Empty, Full;
  wire   \Queue[4][31] , \Queue[4][30] , \Queue[4][29] , \Queue[4][28] ,
         \Queue[4][27] , \Queue[4][26] , \Queue[4][25] , \Queue[4][24] ,
         \Queue[4][23] , \Queue[4][22] , \Queue[4][21] , \Queue[4][20] ,
         \Queue[4][19] , \Queue[4][18] , \Queue[4][17] , \Queue[4][16] ,
         \Queue[4][15] , \Queue[4][14] , \Queue[4][13] , \Queue[4][12] ,
         \Queue[4][11] , \Queue[4][10] , \Queue[4][9] , \Queue[4][8] ,
         \Queue[4][7] , \Queue[4][6] , \Queue[4][5] , \Queue[4][4] ,
         \Queue[4][3] , \Queue[4][2] , \Queue[4][1] , \Queue[4][0] ,
         \Queue[3][31] , \Queue[3][30] , \Queue[3][29] , \Queue[3][28] ,
         \Queue[3][27] , \Queue[3][26] , \Queue[3][25] , \Queue[3][24] ,
         \Queue[3][23] , \Queue[3][22] , \Queue[3][21] , \Queue[3][20] ,
         \Queue[3][19] , \Queue[3][18] , \Queue[3][17] , \Queue[3][16] ,
         \Queue[3][15] , \Queue[3][14] , \Queue[3][13] , \Queue[3][12] ,
         \Queue[3][11] , \Queue[3][10] , \Queue[3][9] , \Queue[3][8] ,
         \Queue[3][7] , \Queue[3][6] , \Queue[3][5] , \Queue[3][4] ,
         \Queue[3][3] , \Queue[3][2] , \Queue[3][1] , \Queue[3][0] ,
         \Queue[2][31] , \Queue[2][30] , \Queue[2][29] , \Queue[2][28] ,
         \Queue[2][27] , \Queue[2][26] , \Queue[2][25] , \Queue[2][24] ,
         \Queue[2][23] , \Queue[2][22] , \Queue[2][21] , \Queue[2][20] ,
         \Queue[2][19] , \Queue[2][18] , \Queue[2][17] , \Queue[2][16] ,
         \Queue[2][15] , \Queue[2][14] , \Queue[2][13] , \Queue[2][12] ,
         \Queue[2][11] , \Queue[2][10] , \Queue[2][9] , \Queue[2][8] ,
         \Queue[2][7] , \Queue[2][6] , \Queue[2][5] , \Queue[2][4] ,
         \Queue[2][3] , \Queue[2][2] , \Queue[2][1] , \Queue[2][0] ,
         \Queue[1][31] , \Queue[1][30] , \Queue[1][29] , \Queue[1][28] ,
         \Queue[1][27] , \Queue[1][26] , \Queue[1][25] , \Queue[1][24] ,
         \Queue[1][23] , \Queue[1][22] , \Queue[1][21] , \Queue[1][20] ,
         \Queue[1][19] , \Queue[1][18] , \Queue[1][17] , \Queue[1][16] ,
         \Queue[1][15] , \Queue[1][14] , \Queue[1][13] , \Queue[1][12] ,
         \Queue[1][11] , \Queue[1][10] , \Queue[1][9] , \Queue[1][8] ,
         \Queue[1][7] , \Queue[1][6] , \Queue[1][5] , \Queue[1][4] ,
         \Queue[1][3] , \Queue[1][2] , \Queue[1][1] , \Queue[1][0] , n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542;
  wire   [2:0] Count;

  FDN2QM1P \Count_reg[0]  ( .D(n377), .CPN(Clk_r), .CD(Rst_n), .Q(Count[0]) );
  FDN2QM1P \Count_reg[1]  ( .D(n378), .CPN(Clk_r), .CD(Rst_n), .Q(Count[1]) );
  FDN2QM1P \Count_reg[2]  ( .D(n379), .CPN(Clk_r), .CD(Rst_n), .Q(Count[2]) );
  FDN1QM1P \Queue_reg[4][30]  ( .D(n411), .CPN(Clk_r), .Q(\Queue[4][30] ) );
  FDN1QM1P \Queue_reg[3][30]  ( .D(n539), .CPN(Clk_r), .Q(\Queue[3][30] ) );
  FDN1QM1P \Queue_reg[2][30]  ( .D(n507), .CPN(Clk_r), .Q(\Queue[2][30] ) );
  FDN1QM1P \Queue_reg[4][29]  ( .D(n410), .CPN(Clk_r), .Q(\Queue[4][29] ) );
  FDN1QM1P \Queue_reg[3][29]  ( .D(n538), .CPN(Clk_r), .Q(\Queue[3][29] ) );
  FDN1QM1P \Queue_reg[2][29]  ( .D(n506), .CPN(Clk_r), .Q(\Queue[2][29] ) );
  FDN1QM1P \Queue_reg[4][28]  ( .D(n409), .CPN(Clk_r), .Q(\Queue[4][28] ) );
  FDN1QM1P \Queue_reg[3][28]  ( .D(n537), .CPN(Clk_r), .Q(\Queue[3][28] ) );
  FDN1QM1P \Queue_reg[2][28]  ( .D(n505), .CPN(Clk_r), .Q(\Queue[2][28] ) );
  FDN1QM1P \Queue_reg[4][27]  ( .D(n408), .CPN(Clk_r), .Q(\Queue[4][27] ) );
  FDN1QM1P \Queue_reg[3][27]  ( .D(n536), .CPN(Clk_r), .Q(\Queue[3][27] ) );
  FDN1QM1P \Queue_reg[2][27]  ( .D(n504), .CPN(Clk_r), .Q(\Queue[2][27] ) );
  FDN1QM1P \Queue_reg[4][26]  ( .D(n407), .CPN(Clk_r), .Q(\Queue[4][26] ) );
  FDN1QM1P \Queue_reg[3][26]  ( .D(n535), .CPN(Clk_r), .Q(\Queue[3][26] ) );
  FDN1QM1P \Queue_reg[2][26]  ( .D(n503), .CPN(Clk_r), .Q(\Queue[2][26] ) );
  FDN1QM1P \Queue_reg[4][25]  ( .D(n406), .CPN(Clk_r), .Q(\Queue[4][25] ) );
  FDN1QM1P \Queue_reg[3][25]  ( .D(n534), .CPN(Clk_r), .Q(\Queue[3][25] ) );
  FDN1QM1P \Queue_reg[2][25]  ( .D(n502), .CPN(Clk_r), .Q(\Queue[2][25] ) );
  FDN1QM1P \Queue_reg[4][24]  ( .D(n405), .CPN(Clk_r), .Q(\Queue[4][24] ) );
  FDN1QM1P \Queue_reg[3][24]  ( .D(n533), .CPN(Clk_r), .Q(\Queue[3][24] ) );
  FDN1QM1P \Queue_reg[2][24]  ( .D(n501), .CPN(Clk_r), .Q(\Queue[2][24] ) );
  FDN1QM1P \Queue_reg[4][23]  ( .D(n404), .CPN(Clk_r), .Q(\Queue[4][23] ) );
  FDN1QM1P \Queue_reg[3][23]  ( .D(n532), .CPN(Clk_r), .Q(\Queue[3][23] ) );
  FDN1QM1P \Queue_reg[2][23]  ( .D(n500), .CPN(Clk_r), .Q(\Queue[2][23] ) );
  FDN1QM1P \Queue_reg[4][22]  ( .D(n403), .CPN(Clk_r), .Q(\Queue[4][22] ) );
  FDN1QM1P \Queue_reg[3][22]  ( .D(n531), .CPN(Clk_r), .Q(\Queue[3][22] ) );
  FDN1QM1P \Queue_reg[2][22]  ( .D(n499), .CPN(Clk_r), .Q(\Queue[2][22] ) );
  FDN1QM1P \Queue_reg[4][21]  ( .D(n402), .CPN(Clk_r), .Q(\Queue[4][21] ) );
  FDN1QM1P \Queue_reg[3][21]  ( .D(n530), .CPN(Clk_r), .Q(\Queue[3][21] ) );
  FDN1QM1P \Queue_reg[2][21]  ( .D(n498), .CPN(Clk_r), .Q(\Queue[2][21] ) );
  FDN1QM1P \Queue_reg[4][20]  ( .D(n401), .CPN(Clk_r), .Q(\Queue[4][20] ) );
  FDN1QM1P \Queue_reg[3][20]  ( .D(n529), .CPN(Clk_r), .Q(\Queue[3][20] ) );
  FDN1QM1P \Queue_reg[2][20]  ( .D(n497), .CPN(Clk_r), .Q(\Queue[2][20] ) );
  FDN1QM1P \Queue_reg[4][19]  ( .D(n400), .CPN(Clk_r), .Q(\Queue[4][19] ) );
  FDN1QM1P \Queue_reg[3][19]  ( .D(n528), .CPN(Clk_r), .Q(\Queue[3][19] ) );
  FDN1QM1P \Queue_reg[2][19]  ( .D(n496), .CPN(Clk_r), .Q(\Queue[2][19] ) );
  FDN1QM1P \Queue_reg[4][18]  ( .D(n399), .CPN(Clk_r), .Q(\Queue[4][18] ) );
  FDN1QM1P \Queue_reg[3][18]  ( .D(n527), .CPN(Clk_r), .Q(\Queue[3][18] ) );
  FDN1QM1P \Queue_reg[2][18]  ( .D(n495), .CPN(Clk_r), .Q(\Queue[2][18] ) );
  FDN1QM1P \Queue_reg[4][17]  ( .D(n398), .CPN(Clk_r), .Q(\Queue[4][17] ) );
  FDN1QM1P \Queue_reg[3][17]  ( .D(n526), .CPN(Clk_r), .Q(\Queue[3][17] ) );
  FDN1QM1P \Queue_reg[2][17]  ( .D(n494), .CPN(Clk_r), .Q(\Queue[2][17] ) );
  FDN1QM1P \Queue_reg[4][16]  ( .D(n397), .CPN(Clk_r), .Q(\Queue[4][16] ) );
  FDN1QM1P \Queue_reg[3][16]  ( .D(n525), .CPN(Clk_r), .Q(\Queue[3][16] ) );
  FDN1QM1P \Queue_reg[2][16]  ( .D(n493), .CPN(Clk_r), .Q(\Queue[2][16] ) );
  FDN1QM1P \Queue_reg[4][15]  ( .D(n396), .CPN(Clk_r), .Q(\Queue[4][15] ) );
  FDN1QM1P \Queue_reg[3][15]  ( .D(n524), .CPN(Clk_r), .Q(\Queue[3][15] ) );
  FDN1QM1P \Queue_reg[2][15]  ( .D(n492), .CPN(Clk_r), .Q(\Queue[2][15] ) );
  FDN1QM1P \Queue_reg[4][14]  ( .D(n395), .CPN(Clk_r), .Q(\Queue[4][14] ) );
  FDN1QM1P \Queue_reg[3][14]  ( .D(n523), .CPN(Clk_r), .Q(\Queue[3][14] ) );
  FDN1QM1P \Queue_reg[2][14]  ( .D(n491), .CPN(Clk_r), .Q(\Queue[2][14] ) );
  FDN1QM1P \Queue_reg[4][13]  ( .D(n394), .CPN(Clk_r), .Q(\Queue[4][13] ) );
  FDN1QM1P \Queue_reg[3][13]  ( .D(n522), .CPN(Clk_r), .Q(\Queue[3][13] ) );
  FDN1QM1P \Queue_reg[2][13]  ( .D(n490), .CPN(Clk_r), .Q(\Queue[2][13] ) );
  FDN1QM1P \Queue_reg[4][12]  ( .D(n393), .CPN(Clk_r), .Q(\Queue[4][12] ) );
  FDN1QM1P \Queue_reg[3][12]  ( .D(n521), .CPN(Clk_r), .Q(\Queue[3][12] ) );
  FDN1QM1P \Queue_reg[2][12]  ( .D(n489), .CPN(Clk_r), .Q(\Queue[2][12] ) );
  FDN1QM1P \Queue_reg[4][11]  ( .D(n392), .CPN(Clk_r), .Q(\Queue[4][11] ) );
  FDN1QM1P \Queue_reg[3][11]  ( .D(n520), .CPN(Clk_r), .Q(\Queue[3][11] ) );
  FDN1QM1P \Queue_reg[2][11]  ( .D(n488), .CPN(Clk_r), .Q(\Queue[2][11] ) );
  FDN1QM1P \Queue_reg[4][10]  ( .D(n391), .CPN(Clk_r), .Q(\Queue[4][10] ) );
  FDN1QM1P \Queue_reg[3][10]  ( .D(n519), .CPN(Clk_r), .Q(\Queue[3][10] ) );
  FDN1QM1P \Queue_reg[2][10]  ( .D(n487), .CPN(Clk_r), .Q(\Queue[2][10] ) );
  FDN1QM1P \Queue_reg[4][9]  ( .D(n390), .CPN(Clk_r), .Q(\Queue[4][9] ) );
  FDN1QM1P \Queue_reg[3][9]  ( .D(n518), .CPN(Clk_r), .Q(\Queue[3][9] ) );
  FDN1QM1P \Queue_reg[2][9]  ( .D(n486), .CPN(Clk_r), .Q(\Queue[2][9] ) );
  FDN1QM1P \Queue_reg[4][8]  ( .D(n389), .CPN(Clk_r), .Q(\Queue[4][8] ) );
  FDN1QM1P \Queue_reg[3][8]  ( .D(n517), .CPN(Clk_r), .Q(\Queue[3][8] ) );
  FDN1QM1P \Queue_reg[2][8]  ( .D(n485), .CPN(Clk_r), .Q(\Queue[2][8] ) );
  FDN1QM1P \Queue_reg[4][7]  ( .D(n388), .CPN(Clk_r), .Q(\Queue[4][7] ) );
  FDN1QM1P \Queue_reg[3][7]  ( .D(n516), .CPN(Clk_r), .Q(\Queue[3][7] ) );
  FDN1QM1P \Queue_reg[2][7]  ( .D(n484), .CPN(Clk_r), .Q(\Queue[2][7] ) );
  FDN1QM1P \Queue_reg[4][6]  ( .D(n387), .CPN(Clk_r), .Q(\Queue[4][6] ) );
  FDN1QM1P \Queue_reg[3][6]  ( .D(n515), .CPN(Clk_r), .Q(\Queue[3][6] ) );
  FDN1QM1P \Queue_reg[2][6]  ( .D(n483), .CPN(Clk_r), .Q(\Queue[2][6] ) );
  FDN1QM1P \Queue_reg[4][5]  ( .D(n386), .CPN(Clk_r), .Q(\Queue[4][5] ) );
  FDN1QM1P \Queue_reg[3][5]  ( .D(n514), .CPN(Clk_r), .Q(\Queue[3][5] ) );
  FDN1QM1P \Queue_reg[2][5]  ( .D(n482), .CPN(Clk_r), .Q(\Queue[2][5] ) );
  FDN1QM1P \Queue_reg[4][4]  ( .D(n385), .CPN(Clk_r), .Q(\Queue[4][4] ) );
  FDN1QM1P \Queue_reg[3][4]  ( .D(n513), .CPN(Clk_r), .Q(\Queue[3][4] ) );
  FDN1QM1P \Queue_reg[2][4]  ( .D(n481), .CPN(Clk_r), .Q(\Queue[2][4] ) );
  FDN1QM1P \Queue_reg[4][3]  ( .D(n384), .CPN(Clk_r), .Q(\Queue[4][3] ) );
  FDN1QM1P \Queue_reg[3][3]  ( .D(n512), .CPN(Clk_r), .Q(\Queue[3][3] ) );
  FDN1QM1P \Queue_reg[2][3]  ( .D(n480), .CPN(Clk_r), .Q(\Queue[2][3] ) );
  FDN1QM1P \Queue_reg[4][2]  ( .D(n383), .CPN(Clk_r), .Q(\Queue[4][2] ) );
  FDN1QM1P \Queue_reg[3][2]  ( .D(n511), .CPN(Clk_r), .Q(\Queue[3][2] ) );
  FDN1QM1P \Queue_reg[2][2]  ( .D(n479), .CPN(Clk_r), .Q(\Queue[2][2] ) );
  FDN1QM1P \Queue_reg[4][1]  ( .D(n382), .CPN(Clk_r), .Q(\Queue[4][1] ) );
  FDN1QM1P \Queue_reg[3][1]  ( .D(n510), .CPN(Clk_r), .Q(\Queue[3][1] ) );
  FDN1QM1P \Queue_reg[2][1]  ( .D(n478), .CPN(Clk_r), .Q(\Queue[2][1] ) );
  FDN1QM1P \Queue_reg[4][0]  ( .D(n381), .CPN(Clk_r), .Q(\Queue[4][0] ) );
  FDN1QM1P \Queue_reg[3][0]  ( .D(n509), .CPN(Clk_r), .Q(\Queue[3][0] ) );
  FDN1QM1P \Queue_reg[2][0]  ( .D(n477), .CPN(Clk_r), .Q(\Queue[2][0] ) );
  FDN1QM1P \Queue_reg[4][31]  ( .D(n380), .CPN(Clk_r), .Q(\Queue[4][31] ) );
  FDN1QM1P \Queue_reg[3][31]  ( .D(n540), .CPN(Clk_r), .Q(\Queue[3][31] ) );
  FDN1QM1P \Queue_reg[2][31]  ( .D(n508), .CPN(Clk_r), .Q(\Queue[2][31] ) );
  FDN2QM1P Full_reg ( .D(n412), .CPN(Clk_r), .CD(Rst_n), .Q(Full) );
  FDN1QM1P \Queue_reg[1][31]  ( .D(n444), .CPN(Clk_r), .Q(\Queue[1][31] ) );
  FDN1QM1P \Queue_reg[0][31]  ( .D(n476), .CPN(Clk_r), .Q(Packet_Out[31]) );
  FDN1QM1P \Queue_reg[1][30]  ( .D(n443), .CPN(Clk_r), .Q(\Queue[1][30] ) );
  FDN1QM1P \Queue_reg[0][30]  ( .D(n475), .CPN(Clk_r), .Q(Packet_Out[30]) );
  FDN1QM1P \Queue_reg[1][29]  ( .D(n442), .CPN(Clk_r), .Q(\Queue[1][29] ) );
  FDN1QM1P \Queue_reg[0][29]  ( .D(n474), .CPN(Clk_r), .Q(Packet_Out[29]) );
  FDN1QM1P \Queue_reg[1][28]  ( .D(n441), .CPN(Clk_r), .Q(\Queue[1][28] ) );
  FDN1QM1P \Queue_reg[0][28]  ( .D(n473), .CPN(Clk_r), .Q(Packet_Out[28]) );
  FDN1QM1P \Queue_reg[1][27]  ( .D(n440), .CPN(Clk_r), .Q(\Queue[1][27] ) );
  FDN1QM1P \Queue_reg[0][27]  ( .D(n472), .CPN(Clk_r), .Q(Packet_Out[27]) );
  FDN1QM1P \Queue_reg[1][26]  ( .D(n439), .CPN(Clk_r), .Q(\Queue[1][26] ) );
  FDN1QM1P \Queue_reg[0][26]  ( .D(n471), .CPN(Clk_r), .Q(Packet_Out[26]) );
  FDN1QM1P \Queue_reg[1][25]  ( .D(n438), .CPN(Clk_r), .Q(\Queue[1][25] ) );
  FDN1QM1P \Queue_reg[0][25]  ( .D(n470), .CPN(Clk_r), .Q(Packet_Out[25]) );
  FDN1QM1P \Queue_reg[1][24]  ( .D(n437), .CPN(Clk_r), .Q(\Queue[1][24] ) );
  FDN1QM1P \Queue_reg[0][24]  ( .D(n469), .CPN(Clk_r), .Q(Packet_Out[24]) );
  FDN1QM1P \Queue_reg[1][23]  ( .D(n436), .CPN(Clk_r), .Q(\Queue[1][23] ) );
  FDN1QM1P \Queue_reg[0][23]  ( .D(n468), .CPN(Clk_r), .Q(Packet_Out[23]) );
  FDN1QM1P \Queue_reg[1][22]  ( .D(n435), .CPN(Clk_r), .Q(\Queue[1][22] ) );
  FDN1QM1P \Queue_reg[0][22]  ( .D(n467), .CPN(Clk_r), .Q(Packet_Out[22]) );
  FDN1QM1P \Queue_reg[1][21]  ( .D(n434), .CPN(Clk_r), .Q(\Queue[1][21] ) );
  FDN1QM1P \Queue_reg[0][21]  ( .D(n466), .CPN(Clk_r), .Q(Packet_Out[21]) );
  FDN1QM1P \Queue_reg[1][20]  ( .D(n433), .CPN(Clk_r), .Q(\Queue[1][20] ) );
  FDN1QM1P \Queue_reg[0][20]  ( .D(n465), .CPN(Clk_r), .Q(Packet_Out[20]) );
  FDN1QM1P \Queue_reg[1][19]  ( .D(n432), .CPN(Clk_r), .Q(\Queue[1][19] ) );
  FDN1QM1P \Queue_reg[0][19]  ( .D(n464), .CPN(Clk_r), .Q(Packet_Out[19]) );
  FDN1QM1P \Queue_reg[1][18]  ( .D(n431), .CPN(Clk_r), .Q(\Queue[1][18] ) );
  FDN1QM1P \Queue_reg[0][18]  ( .D(n463), .CPN(Clk_r), .Q(Packet_Out[18]) );
  FDN1QM1P \Queue_reg[1][17]  ( .D(n430), .CPN(Clk_r), .Q(\Queue[1][17] ) );
  FDN1QM1P \Queue_reg[0][17]  ( .D(n462), .CPN(Clk_r), .Q(Packet_Out[17]) );
  FDN1QM1P \Queue_reg[1][16]  ( .D(n429), .CPN(Clk_r), .Q(\Queue[1][16] ) );
  FDN1QM1P \Queue_reg[0][16]  ( .D(n461), .CPN(Clk_r), .Q(Packet_Out[16]) );
  FDN1QM1P \Queue_reg[1][15]  ( .D(n428), .CPN(Clk_r), .Q(\Queue[1][15] ) );
  FDN1QM1P \Queue_reg[0][15]  ( .D(n460), .CPN(Clk_r), .Q(Packet_Out[15]) );
  FDN1QM1P \Queue_reg[1][14]  ( .D(n427), .CPN(Clk_r), .Q(\Queue[1][14] ) );
  FDN1QM1P \Queue_reg[0][14]  ( .D(n459), .CPN(Clk_r), .Q(Packet_Out[14]) );
  FDN1QM1P \Queue_reg[1][13]  ( .D(n426), .CPN(Clk_r), .Q(\Queue[1][13] ) );
  FDN1QM1P \Queue_reg[0][13]  ( .D(n458), .CPN(Clk_r), .Q(Packet_Out[13]) );
  FDN1QM1P \Queue_reg[1][12]  ( .D(n425), .CPN(Clk_r), .Q(\Queue[1][12] ) );
  FDN1QM1P \Queue_reg[0][12]  ( .D(n457), .CPN(Clk_r), .Q(Packet_Out[12]) );
  FDN1QM1P \Queue_reg[1][11]  ( .D(n424), .CPN(Clk_r), .Q(\Queue[1][11] ) );
  FDN1QM1P \Queue_reg[0][11]  ( .D(n456), .CPN(Clk_r), .Q(Packet_Out[11]) );
  FDN1QM1P \Queue_reg[1][10]  ( .D(n423), .CPN(Clk_r), .Q(\Queue[1][10] ) );
  FDN1QM1P \Queue_reg[0][10]  ( .D(n455), .CPN(Clk_r), .Q(Packet_Out[10]) );
  FDN1QM1P \Queue_reg[1][9]  ( .D(n422), .CPN(Clk_r), .Q(\Queue[1][9] ) );
  FDN1QM1P \Queue_reg[0][9]  ( .D(n454), .CPN(Clk_r), .Q(Packet_Out[9]) );
  FDN1QM1P \Queue_reg[1][8]  ( .D(n421), .CPN(Clk_r), .Q(\Queue[1][8] ) );
  FDN1QM1P \Queue_reg[0][8]  ( .D(n453), .CPN(Clk_r), .Q(Packet_Out[8]) );
  FDN1QM1P \Queue_reg[1][7]  ( .D(n420), .CPN(Clk_r), .Q(\Queue[1][7] ) );
  FDN1QM1P \Queue_reg[0][7]  ( .D(n452), .CPN(Clk_r), .Q(Packet_Out[7]) );
  FDN1QM1P \Queue_reg[1][6]  ( .D(n419), .CPN(Clk_r), .Q(\Queue[1][6] ) );
  FDN1QM1P \Queue_reg[0][6]  ( .D(n451), .CPN(Clk_r), .Q(Packet_Out[6]) );
  FDN1QM1P \Queue_reg[1][5]  ( .D(n418), .CPN(Clk_r), .Q(\Queue[1][5] ) );
  FDN1QM1P \Queue_reg[0][5]  ( .D(n450), .CPN(Clk_r), .Q(Packet_Out[5]) );
  FDN1QM1P \Queue_reg[1][4]  ( .D(n417), .CPN(Clk_r), .Q(\Queue[1][4] ) );
  FDN1QM1P \Queue_reg[0][4]  ( .D(n449), .CPN(Clk_r), .Q(Packet_Out[4]) );
  FDN1QM1P \Queue_reg[1][3]  ( .D(n416), .CPN(Clk_r), .Q(\Queue[1][3] ) );
  FDN1QM1P \Queue_reg[0][3]  ( .D(n448), .CPN(Clk_r), .Q(Packet_Out[3]) );
  FDN1QM1P \Queue_reg[1][2]  ( .D(n415), .CPN(Clk_r), .Q(\Queue[1][2] ) );
  FDN1QM1P \Queue_reg[0][2]  ( .D(n447), .CPN(Clk_r), .Q(Packet_Out[2]) );
  FDN1QM1P \Queue_reg[1][1]  ( .D(n414), .CPN(Clk_r), .Q(\Queue[1][1] ) );
  FDN1QM1P \Queue_reg[0][1]  ( .D(n446), .CPN(Clk_r), .Q(Packet_Out[1]) );
  FDN1QM1P \Queue_reg[1][0]  ( .D(n413), .CPN(Clk_r), .Q(\Queue[1][0] ) );
  FDN1QM1P \Queue_reg[0][0]  ( .D(n445), .CPN(Clk_r), .Q(Packet_Out[0]) );
  FDN2QM1P Empty_reg ( .D(n542), .CPN(Clk_r), .CD(Rst_n), .Q(n541) );
  NR3M1P U3 ( .A(Count[0]), .B(Count[2]), .C(n22), .Z(n100) );
  BUFM2P U4 ( .A(n97), .Z(n9) );
  BUFM1P U5 ( .A(n97), .Z(n10) );
  BUFM1P U6 ( .A(n205), .Z(n12) );
  BUFM2P U7 ( .A(n132), .Z(n3) );
  BUFM1P U8 ( .A(n205), .Z(n11) );
  NR3M1P U9 ( .A(n23), .B(Count[2]), .C(Count[1]), .Z(n376) );
  N1M1P U10 ( .A(Read_Ack), .Z(n137) );
  NR3M1P U11 ( .A(Count[2]), .B(n23), .C(n22), .Z(n140) );
  N1M1P U12 ( .A(n4), .Z(n99) );
  AOI21M2P U13 ( .A(n4), .B(n376), .C(n141), .Z(n95) );
  AOI21M3P U14 ( .A(n4), .B(n100), .C(n141), .Z(n57) );
  OAI211M4P U15 ( .A(n100), .B(n137), .C(n4), .D(n24), .Z(n59) );
  NR2FM3P U16 ( .A(n61), .B(n21), .Z(n20) );
  OAI211M4P U17 ( .A(n142), .B(n137), .C(n4), .D(n136), .Z(n208) );
  OAI211M4P U18 ( .A(n140), .B(n137), .C(n4), .D(n98), .Z(n135) );
  OAI21M2P U19 ( .A(n4), .B(Read_Ack), .C(n24), .Z(n56) );
  N1M1P U20 ( .A(n142), .Z(n21) );
  NR3M1P U21 ( .A(Count[0]), .B(Count[1]), .C(n19), .Z(n142) );
  N1M1P U22 ( .A(Count[2]), .Z(n19) );
  N1M1P U23 ( .A(Count[0]), .Z(n23) );
  N1M1P U24 ( .A(Count[1]), .Z(n22) );
  BUFM2P U25 ( .A(n95), .Z(n8) );
  AOI21M6P U26 ( .A(n4), .B(n142), .C(n141), .Z(n205) );
  ND2M2P U27 ( .A(Read_Ack), .B(Rst_n), .Z(n141) );
  ND2M2P U28 ( .A(n18), .B(Rst_n), .Z(n61) );
  NR2M3P U29 ( .A(Read_Ack), .B(n99), .Z(n18) );
  BUFM10P U30 ( .A(Write_Ack), .Z(n4) );
  OAI211M4P U31 ( .A(n100), .B(n139), .C(Rst_n), .D(n138), .Z(n133) );
  N1M1P U32 ( .A(Packet_In[23]), .Z(n190) );
  N1M1P U33 ( .A(Packet_In[25]), .Z(n194) );
  N1M1P U34 ( .A(Packet_In[28]), .Z(n200) );
  N1M1P U35 ( .A(Packet_In[27]), .Z(n198) );
  N1M1P U36 ( .A(Packet_In[26]), .Z(n196) );
  N1M1P U37 ( .A(Packet_In[29]), .Z(n202) );
  OAI211M4P U38 ( .A(n140), .B(n139), .C(Rst_n), .D(n138), .Z(n206) );
  N1M1P U39 ( .A(Packet_In[31]), .Z(n373) );
  N1M1P U40 ( .A(Packet_In[24]), .Z(n192) );
  N1M1P U41 ( .A(Packet_In[20]), .Z(n184) );
  N1M1P U42 ( .A(Packet_In[21]), .Z(n186) );
  N1M1P U43 ( .A(Packet_In[22]), .Z(n188) );
  N1M1P U44 ( .A(Packet_In[0]), .Z(n144) );
  N1M1P U45 ( .A(Packet_In[12]), .Z(n168) );
  N1M1P U46 ( .A(Packet_In[3]), .Z(n150) );
  N1M1P U47 ( .A(Packet_In[4]), .Z(n152) );
  N1M1P U48 ( .A(Packet_In[5]), .Z(n154) );
  N1M1P U49 ( .A(Packet_In[14]), .Z(n172) );
  N1M1P U50 ( .A(Packet_In[6]), .Z(n156) );
  N1M1P U51 ( .A(Packet_In[30]), .Z(n204) );
  N1M1P U52 ( .A(Packet_In[17]), .Z(n178) );
  N1M1P U53 ( .A(Packet_In[1]), .Z(n146) );
  N1M1P U54 ( .A(Packet_In[2]), .Z(n148) );
  N1M1P U55 ( .A(Packet_In[7]), .Z(n158) );
  N1M1P U56 ( .A(Packet_In[9]), .Z(n162) );
  N1M1P U57 ( .A(Packet_In[19]), .Z(n182) );
  N1M1P U58 ( .A(Packet_In[15]), .Z(n174) );
  N1M1P U59 ( .A(Packet_In[8]), .Z(n160) );
  N1M1P U60 ( .A(Packet_In[13]), .Z(n170) );
  N1M1P U61 ( .A(Packet_In[16]), .Z(n176) );
  N1M1P U62 ( .A(Packet_In[11]), .Z(n166) );
  N1M1P U63 ( .A(Packet_In[10]), .Z(n164) );
  N1M1P U64 ( .A(Packet_In[18]), .Z(n180) );
  BUFM2P U65 ( .A(n57), .Z(n7) );
  BUFM2P U66 ( .A(n56), .Z(n6) );
  BUFM2P U67 ( .A(n56), .Z(n5) );
  N1M2P U68 ( .A(n18), .Z(n139) );
  N1M2P U69 ( .A(n62), .Z(n94) );
  OAI211M1P U70 ( .A(n376), .B(n137), .C(n4), .D(n62), .Z(n97) );
  NR2M1P U71 ( .A(n137), .B(n4), .Z(n375) );
  NR2M1P U72 ( .A(n18), .B(n375), .Z(n374) );
  AOI22CDNM1P U73 ( .A(n374), .B(n23), .C(n374), .D(n23), .Z(n377) );
  N1M1P U74 ( .A(n375), .Z(n17) );
  AOI22M1P U75 ( .A(Count[0]), .B(n139), .C(n17), .D(n23), .Z(n14) );
  AOI22CDNM1P U76 ( .A(Count[1]), .B(n14), .C(n14), .D(Count[1]), .Z(n378) );
  ND3M1P U77 ( .A(n23), .B(n19), .C(n22), .Z(n60) );
  ND2M1P U78 ( .A(Count[1]), .B(Read_Ack), .Z(n13) );
  OAI211M1P U79 ( .A(Count[1]), .B(n139), .C(n14), .D(n13), .Z(n15) );
  AOI22M1P U80 ( .A(n18), .B(n140), .C(Count[2]), .D(n15), .Z(n16) );
  OAI21M1P U81 ( .A(n60), .B(n17), .C(n16), .Z(n379) );
  AOI22CDNM1P U82 ( .A(n20), .B(n373), .C(\Queue[4][31] ), .D(n20), .Z(n380)
         );
  AOI22CDNM1P U83 ( .A(n20), .B(n144), .C(\Queue[4][0] ), .D(n20), .Z(n381) );
  AOI22CDNM1P U84 ( .A(n20), .B(n146), .C(\Queue[4][1] ), .D(n20), .Z(n382) );
  AOI22CDNM1P U85 ( .A(n20), .B(n148), .C(\Queue[4][2] ), .D(n20), .Z(n383) );
  AOI22CDNM1P U86 ( .A(n20), .B(n150), .C(\Queue[4][3] ), .D(n20), .Z(n384) );
  AOI22CDNM1P U87 ( .A(n20), .B(n152), .C(\Queue[4][4] ), .D(n20), .Z(n385) );
  AOI22CDNM1P U88 ( .A(n20), .B(n154), .C(\Queue[4][5] ), .D(n20), .Z(n386) );
  AOI22CDNM1P U89 ( .A(n20), .B(n156), .C(\Queue[4][6] ), .D(n20), .Z(n387) );
  AOI22CDNM1P U90 ( .A(n20), .B(n158), .C(\Queue[4][7] ), .D(n20), .Z(n388) );
  AOI22CDNM1P U91 ( .A(n20), .B(n160), .C(\Queue[4][8] ), .D(n20), .Z(n389) );
  AOI22CDNM1P U92 ( .A(n20), .B(n162), .C(\Queue[4][9] ), .D(n20), .Z(n390) );
  AOI22CDNM1P U93 ( .A(n20), .B(n164), .C(\Queue[4][10] ), .D(n20), .Z(n391)
         );
  AOI22CDNM1P U94 ( .A(n20), .B(n166), .C(\Queue[4][11] ), .D(n20), .Z(n392)
         );
  AOI22CDNM1P U95 ( .A(n20), .B(n168), .C(\Queue[4][12] ), .D(n20), .Z(n393)
         );
  AOI22CDNM1P U96 ( .A(n20), .B(n170), .C(\Queue[4][13] ), .D(n20), .Z(n394)
         );
  AOI22CDNM1P U97 ( .A(n20), .B(n172), .C(\Queue[4][14] ), .D(n20), .Z(n395)
         );
  AOI22CDNM1P U98 ( .A(n20), .B(n174), .C(\Queue[4][15] ), .D(n20), .Z(n396)
         );
  AOI22CDNM1P U99 ( .A(n20), .B(n176), .C(\Queue[4][16] ), .D(n20), .Z(n397)
         );
  AOI22CDNM1P U100 ( .A(n20), .B(n178), .C(\Queue[4][17] ), .D(n20), .Z(n398)
         );
  AOI22CDNM1P U101 ( .A(n20), .B(n180), .C(\Queue[4][18] ), .D(n20), .Z(n399)
         );
  AOI22CDNM1P U102 ( .A(n20), .B(n182), .C(\Queue[4][19] ), .D(n20), .Z(n400)
         );
  AOI22CDNM1P U103 ( .A(n20), .B(n184), .C(\Queue[4][20] ), .D(n20), .Z(n401)
         );
  AOI22CDNM1P U104 ( .A(n20), .B(n186), .C(\Queue[4][21] ), .D(n20), .Z(n402)
         );
  AOI22CDNM1P U105 ( .A(n20), .B(n188), .C(\Queue[4][22] ), .D(n20), .Z(n403)
         );
  AOI22CDNM1P U106 ( .A(n20), .B(n190), .C(\Queue[4][23] ), .D(n20), .Z(n404)
         );
  AOI22CDNM1P U107 ( .A(n20), .B(n192), .C(\Queue[4][24] ), .D(n20), .Z(n405)
         );
  AOI22CDNM1P U108 ( .A(n20), .B(n194), .C(\Queue[4][25] ), .D(n20), .Z(n406)
         );
  AOI22CDNM1P U109 ( .A(n20), .B(n196), .C(\Queue[4][26] ), .D(n20), .Z(n407)
         );
  AOI22CDNM1P U110 ( .A(n20), .B(n198), .C(\Queue[4][27] ), .D(n20), .Z(n408)
         );
  AOI22CDNM1P U111 ( .A(n20), .B(n200), .C(\Queue[4][28] ), .D(n20), .Z(n409)
         );
  AOI22CDNM1P U112 ( .A(n20), .B(n202), .C(\Queue[4][29] ), .D(n20), .Z(n410)
         );
  AOI22CDNM1P U113 ( .A(n20), .B(n204), .C(\Queue[4][30] ), .D(n20), .Z(n411)
         );
  OAI22CDNM1P U114 ( .A(n139), .B(n21), .C(n374), .D(Full), .Z(n412) );
  OA21M1P U115 ( .A(n139), .B(n376), .C(Rst_n), .Z(n24) );
  AOI22M1P U116 ( .A(\Queue[2][0] ), .B(n57), .C(\Queue[1][0] ), .D(n5), .Z(
        n25) );
  OAI21M1P U117 ( .A(n144), .B(n59), .C(n25), .Z(n413) );
  AOI22M1P U118 ( .A(n7), .B(\Queue[2][1] ), .C(\Queue[1][1] ), .D(n5), .Z(n26) );
  OAI21M1P U119 ( .A(n59), .B(n146), .C(n26), .Z(n414) );
  AOI22M1P U120 ( .A(n57), .B(\Queue[2][2] ), .C(\Queue[1][2] ), .D(n5), .Z(
        n27) );
  OAI21M1P U121 ( .A(n59), .B(n148), .C(n27), .Z(n415) );
  AOI22M1P U122 ( .A(n57), .B(\Queue[2][3] ), .C(\Queue[1][3] ), .D(n5), .Z(
        n28) );
  OAI21M1P U123 ( .A(n59), .B(n150), .C(n28), .Z(n416) );
  AOI22M1P U124 ( .A(n57), .B(\Queue[2][4] ), .C(\Queue[1][4] ), .D(n5), .Z(
        n29) );
  OAI21M1P U125 ( .A(n59), .B(n152), .C(n29), .Z(n417) );
  AOI22M1P U126 ( .A(n57), .B(\Queue[2][5] ), .C(\Queue[1][5] ), .D(n5), .Z(
        n30) );
  OAI21M1P U127 ( .A(n59), .B(n154), .C(n30), .Z(n418) );
  AOI22M1P U128 ( .A(n57), .B(\Queue[2][6] ), .C(\Queue[1][6] ), .D(n5), .Z(
        n31) );
  OAI21M1P U129 ( .A(n59), .B(n156), .C(n31), .Z(n419) );
  AOI22M1P U130 ( .A(n57), .B(\Queue[2][7] ), .C(\Queue[1][7] ), .D(n5), .Z(
        n32) );
  OAI21M1P U131 ( .A(n59), .B(n158), .C(n32), .Z(n420) );
  AOI22M1P U132 ( .A(n57), .B(\Queue[2][8] ), .C(\Queue[1][8] ), .D(n5), .Z(
        n33) );
  OAI21M1P U133 ( .A(n59), .B(n160), .C(n33), .Z(n421) );
  AOI22M1P U134 ( .A(n7), .B(\Queue[2][9] ), .C(\Queue[1][9] ), .D(n56), .Z(
        n34) );
  OAI21M1P U135 ( .A(n59), .B(n162), .C(n34), .Z(n422) );
  AOI22M1P U136 ( .A(n57), .B(\Queue[2][10] ), .C(\Queue[1][10] ), .D(n5), .Z(
        n35) );
  OAI21M1P U137 ( .A(n59), .B(n164), .C(n35), .Z(n423) );
  AOI22M1P U138 ( .A(n57), .B(\Queue[2][11] ), .C(\Queue[1][11] ), .D(n6), .Z(
        n36) );
  OAI21M1P U139 ( .A(n59), .B(n166), .C(n36), .Z(n424) );
  AOI22M1P U140 ( .A(n7), .B(\Queue[2][12] ), .C(\Queue[1][12] ), .D(n56), .Z(
        n37) );
  OAI21M1P U141 ( .A(n59), .B(n168), .C(n37), .Z(n425) );
  AOI22M1P U142 ( .A(n7), .B(\Queue[2][13] ), .C(\Queue[1][13] ), .D(n56), .Z(
        n38) );
  OAI21M1P U143 ( .A(n59), .B(n170), .C(n38), .Z(n426) );
  AOI22M1P U144 ( .A(n7), .B(\Queue[2][14] ), .C(\Queue[1][14] ), .D(n56), .Z(
        n39) );
  OAI21M1P U145 ( .A(n59), .B(n172), .C(n39), .Z(n427) );
  AOI22M1P U146 ( .A(n7), .B(\Queue[2][15] ), .C(\Queue[1][15] ), .D(n56), .Z(
        n40) );
  OAI21M1P U147 ( .A(n59), .B(n174), .C(n40), .Z(n428) );
  AOI22M1P U148 ( .A(n7), .B(\Queue[2][16] ), .C(\Queue[1][16] ), .D(n56), .Z(
        n41) );
  OAI21M1P U149 ( .A(n59), .B(n176), .C(n41), .Z(n429) );
  AOI22M1P U150 ( .A(n7), .B(\Queue[2][17] ), .C(\Queue[1][17] ), .D(n56), .Z(
        n42) );
  OAI21M1P U151 ( .A(n59), .B(n178), .C(n42), .Z(n430) );
  AOI22M1P U152 ( .A(n7), .B(\Queue[2][18] ), .C(\Queue[1][18] ), .D(n6), .Z(
        n43) );
  OAI21M1P U153 ( .A(n59), .B(n180), .C(n43), .Z(n431) );
  AOI22M1P U154 ( .A(n7), .B(\Queue[2][19] ), .C(\Queue[1][19] ), .D(n6), .Z(
        n44) );
  OAI21M1P U155 ( .A(n59), .B(n182), .C(n44), .Z(n432) );
  AOI22M1P U156 ( .A(n7), .B(\Queue[2][20] ), .C(\Queue[1][20] ), .D(n6), .Z(
        n45) );
  OAI21M1P U157 ( .A(n59), .B(n184), .C(n45), .Z(n433) );
  AOI22M1P U158 ( .A(n7), .B(\Queue[2][21] ), .C(\Queue[1][21] ), .D(n6), .Z(
        n46) );
  OAI21M1P U159 ( .A(n59), .B(n186), .C(n46), .Z(n434) );
  AOI22M1P U160 ( .A(n57), .B(\Queue[2][22] ), .C(\Queue[1][22] ), .D(n6), .Z(
        n47) );
  OAI21M1P U161 ( .A(n59), .B(n188), .C(n47), .Z(n435) );
  AOI22M1P U162 ( .A(n7), .B(\Queue[2][23] ), .C(\Queue[1][23] ), .D(n6), .Z(
        n48) );
  OAI21M1P U163 ( .A(n59), .B(n190), .C(n48), .Z(n436) );
  AOI22M1P U164 ( .A(n57), .B(\Queue[2][24] ), .C(\Queue[1][24] ), .D(n6), .Z(
        n49) );
  OAI21M1P U165 ( .A(n59), .B(n192), .C(n49), .Z(n437) );
  AOI22M1P U166 ( .A(n57), .B(\Queue[2][25] ), .C(\Queue[1][25] ), .D(n6), .Z(
        n50) );
  OAI21M1P U167 ( .A(n59), .B(n194), .C(n50), .Z(n438) );
  AOI22M1P U168 ( .A(n57), .B(\Queue[2][26] ), .C(\Queue[1][26] ), .D(n6), .Z(
        n51) );
  OAI21M1P U169 ( .A(n59), .B(n196), .C(n51), .Z(n439) );
  AOI22M1P U170 ( .A(n57), .B(\Queue[2][27] ), .C(\Queue[1][27] ), .D(n6), .Z(
        n52) );
  OAI21M1P U171 ( .A(n59), .B(n198), .C(n52), .Z(n440) );
  AOI22M1P U172 ( .A(n57), .B(\Queue[2][28] ), .C(\Queue[1][28] ), .D(n5), .Z(
        n53) );
  OAI21M1P U173 ( .A(n59), .B(n200), .C(n53), .Z(n441) );
  AOI22M1P U174 ( .A(n57), .B(\Queue[2][29] ), .C(\Queue[1][29] ), .D(n5), .Z(
        n54) );
  OAI21M1P U175 ( .A(n59), .B(n202), .C(n54), .Z(n442) );
  AOI22M1P U176 ( .A(n57), .B(\Queue[2][30] ), .C(\Queue[1][30] ), .D(n6), .Z(
        n55) );
  OAI21M1P U177 ( .A(n59), .B(n204), .C(n55), .Z(n443) );
  AOI22M1P U178 ( .A(n57), .B(\Queue[2][31] ), .C(\Queue[1][31] ), .D(n5), .Z(
        n58) );
  OAI21M1P U179 ( .A(n59), .B(n373), .C(n58), .Z(n444) );
  OAI21M1P U180 ( .A(n61), .B(n60), .C(n141), .Z(n62) );
  AOI22M1P U181 ( .A(\Queue[1][0] ), .B(n8), .C(n94), .D(Packet_Out[0]), .Z(
        n63) );
  OAI21M1P U182 ( .A(n144), .B(n9), .C(n63), .Z(n445) );
  AOI22M1P U183 ( .A(\Queue[1][1] ), .B(n8), .C(n94), .D(Packet_Out[1]), .Z(
        n64) );
  OAI21M1P U184 ( .A(n146), .B(n9), .C(n64), .Z(n446) );
  AOI22M1P U185 ( .A(\Queue[1][2] ), .B(n8), .C(n94), .D(Packet_Out[2]), .Z(
        n65) );
  OAI21M1P U186 ( .A(n148), .B(n9), .C(n65), .Z(n447) );
  AOI22M1P U187 ( .A(\Queue[1][3] ), .B(n95), .C(n94), .D(Packet_Out[3]), .Z(
        n66) );
  OAI21M1P U188 ( .A(n150), .B(n9), .C(n66), .Z(n448) );
  AOI22M1P U189 ( .A(\Queue[1][4] ), .B(n95), .C(n94), .D(Packet_Out[4]), .Z(
        n67) );
  OAI21M1P U190 ( .A(n152), .B(n9), .C(n67), .Z(n449) );
  AOI22M1P U191 ( .A(\Queue[1][5] ), .B(n95), .C(n94), .D(Packet_Out[5]), .Z(
        n68) );
  OAI21M1P U192 ( .A(n154), .B(n9), .C(n68), .Z(n450) );
  AOI22M1P U193 ( .A(\Queue[1][6] ), .B(n95), .C(n94), .D(Packet_Out[6]), .Z(
        n69) );
  OAI21M1P U194 ( .A(n156), .B(n9), .C(n69), .Z(n451) );
  AOI22M1P U195 ( .A(\Queue[1][7] ), .B(n95), .C(n94), .D(Packet_Out[7]), .Z(
        n70) );
  OAI21M1P U196 ( .A(n158), .B(n9), .C(n70), .Z(n452) );
  AOI22M1P U197 ( .A(\Queue[1][8] ), .B(n95), .C(n94), .D(Packet_Out[8]), .Z(
        n71) );
  OAI21M1P U198 ( .A(n160), .B(n9), .C(n71), .Z(n453) );
  AOI22M1P U199 ( .A(\Queue[1][9] ), .B(n95), .C(n94), .D(Packet_Out[9]), .Z(
        n72) );
  OAI21M1P U200 ( .A(n162), .B(n9), .C(n72), .Z(n454) );
  AOI22M1P U201 ( .A(\Queue[1][10] ), .B(n8), .C(n94), .D(Packet_Out[10]), .Z(
        n73) );
  OAI21M1P U202 ( .A(n164), .B(n9), .C(n73), .Z(n455) );
  AOI22M1P U203 ( .A(\Queue[1][11] ), .B(n8), .C(n94), .D(Packet_Out[11]), .Z(
        n74) );
  OAI21M1P U204 ( .A(n166), .B(n9), .C(n74), .Z(n456) );
  AOI22M1P U205 ( .A(\Queue[1][12] ), .B(n8), .C(n94), .D(Packet_Out[12]), .Z(
        n75) );
  OAI21M1P U206 ( .A(n168), .B(n9), .C(n75), .Z(n457) );
  AOI22M1P U207 ( .A(\Queue[1][13] ), .B(n8), .C(n94), .D(Packet_Out[13]), .Z(
        n76) );
  OAI21M1P U208 ( .A(n170), .B(n9), .C(n76), .Z(n458) );
  AOI22M1P U209 ( .A(\Queue[1][14] ), .B(n8), .C(n94), .D(Packet_Out[14]), .Z(
        n77) );
  OAI21M1P U210 ( .A(n172), .B(n9), .C(n77), .Z(n459) );
  AOI22M1P U211 ( .A(\Queue[1][15] ), .B(n8), .C(n94), .D(Packet_Out[15]), .Z(
        n78) );
  OAI21M1P U212 ( .A(n174), .B(n9), .C(n78), .Z(n460) );
  AOI22M1P U213 ( .A(\Queue[1][16] ), .B(n95), .C(n94), .D(Packet_Out[16]), 
        .Z(n79) );
  OAI21M1P U214 ( .A(n176), .B(n9), .C(n79), .Z(n461) );
  AOI22M1P U215 ( .A(\Queue[1][17] ), .B(n95), .C(n94), .D(Packet_Out[17]), 
        .Z(n80) );
  OAI21M1P U216 ( .A(n178), .B(n9), .C(n80), .Z(n462) );
  AOI22M1P U217 ( .A(\Queue[1][18] ), .B(n95), .C(n94), .D(Packet_Out[18]), 
        .Z(n81) );
  OAI21M1P U218 ( .A(n180), .B(n9), .C(n81), .Z(n463) );
  AOI22M1P U219 ( .A(\Queue[1][19] ), .B(n95), .C(n94), .D(Packet_Out[19]), 
        .Z(n82) );
  OAI21M1P U220 ( .A(n182), .B(n9), .C(n82), .Z(n464) );
  AOI22M1P U221 ( .A(\Queue[1][20] ), .B(n8), .C(n94), .D(Packet_Out[20]), .Z(
        n83) );
  OAI21M1P U222 ( .A(n184), .B(n10), .C(n83), .Z(n465) );
  AOI22M1P U223 ( .A(\Queue[1][21] ), .B(n8), .C(n94), .D(Packet_Out[21]), .Z(
        n84) );
  OAI21M1P U224 ( .A(n186), .B(n10), .C(n84), .Z(n466) );
  AOI22M1P U225 ( .A(\Queue[1][22] ), .B(n8), .C(n94), .D(Packet_Out[22]), .Z(
        n85) );
  OAI21M1P U226 ( .A(n188), .B(n10), .C(n85), .Z(n467) );
  AOI22M1P U227 ( .A(\Queue[1][23] ), .B(n8), .C(n94), .D(Packet_Out[23]), .Z(
        n86) );
  OAI21M1P U228 ( .A(n190), .B(n10), .C(n86), .Z(n468) );
  AOI22M1P U229 ( .A(\Queue[1][24] ), .B(n8), .C(n94), .D(Packet_Out[24]), .Z(
        n87) );
  OAI21M1P U230 ( .A(n192), .B(n10), .C(n87), .Z(n469) );
  AOI22M1P U231 ( .A(\Queue[1][25] ), .B(n8), .C(n94), .D(Packet_Out[25]), .Z(
        n88) );
  OAI21M1P U232 ( .A(n194), .B(n10), .C(n88), .Z(n470) );
  AOI22M1P U233 ( .A(\Queue[1][26] ), .B(n8), .C(n94), .D(Packet_Out[26]), .Z(
        n89) );
  OAI21M1P U234 ( .A(n196), .B(n10), .C(n89), .Z(n471) );
  AOI22M1P U235 ( .A(\Queue[1][27] ), .B(n8), .C(n94), .D(Packet_Out[27]), .Z(
        n90) );
  OAI21M1P U236 ( .A(n198), .B(n10), .C(n90), .Z(n472) );
  AOI22M1P U237 ( .A(\Queue[1][28] ), .B(n8), .C(n94), .D(Packet_Out[28]), .Z(
        n91) );
  OAI21M1P U238 ( .A(n200), .B(n10), .C(n91), .Z(n473) );
  AOI22M1P U239 ( .A(\Queue[1][29] ), .B(n8), .C(n94), .D(Packet_Out[29]), .Z(
        n92) );
  OAI21M1P U240 ( .A(n202), .B(n10), .C(n92), .Z(n474) );
  AOI22M1P U241 ( .A(\Queue[1][30] ), .B(n95), .C(n94), .D(Packet_Out[30]), 
        .Z(n93) );
  OAI21M1P U242 ( .A(n204), .B(n9), .C(n93), .Z(n475) );
  AOI22M1P U243 ( .A(\Queue[1][31] ), .B(n8), .C(n94), .D(Packet_Out[31]), .Z(
        n96) );
  OAI21M1P U244 ( .A(n373), .B(n10), .C(n96), .Z(n476) );
  OA21M1P U245 ( .A(n139), .B(n100), .C(Rst_n), .Z(n98) );
  ND2M1P U246 ( .A(n99), .B(n137), .Z(n138) );
  AOI21M1P U247 ( .A(n4), .B(n140), .C(n141), .Z(n132) );
  AOI22M1P U248 ( .A(\Queue[2][0] ), .B(n133), .C(\Queue[3][0] ), .D(n3), .Z(
        n101) );
  OAI21M1P U249 ( .A(n144), .B(n135), .C(n101), .Z(n477) );
  AOI22M1P U250 ( .A(\Queue[2][1] ), .B(n133), .C(n3), .D(\Queue[3][1] ), .Z(
        n102) );
  OAI21M1P U251 ( .A(n146), .B(n135), .C(n102), .Z(n478) );
  AOI22M1P U252 ( .A(\Queue[2][2] ), .B(n133), .C(n3), .D(\Queue[3][2] ), .Z(
        n103) );
  OAI21M1P U253 ( .A(n148), .B(n135), .C(n103), .Z(n479) );
  AOI22M1P U254 ( .A(\Queue[2][3] ), .B(n133), .C(n3), .D(\Queue[3][3] ), .Z(
        n104) );
  OAI21M1P U255 ( .A(n150), .B(n135), .C(n104), .Z(n480) );
  AOI22M1P U256 ( .A(\Queue[2][4] ), .B(n133), .C(n3), .D(\Queue[3][4] ), .Z(
        n105) );
  OAI21M1P U257 ( .A(n152), .B(n135), .C(n105), .Z(n481) );
  AOI22M1P U258 ( .A(\Queue[2][5] ), .B(n133), .C(n3), .D(\Queue[3][5] ), .Z(
        n106) );
  OAI21M1P U259 ( .A(n154), .B(n135), .C(n106), .Z(n482) );
  AOI22M1P U260 ( .A(\Queue[2][6] ), .B(n133), .C(n3), .D(\Queue[3][6] ), .Z(
        n107) );
  OAI21M1P U261 ( .A(n156), .B(n135), .C(n107), .Z(n483) );
  AOI22M1P U262 ( .A(\Queue[2][7] ), .B(n133), .C(n3), .D(\Queue[3][7] ), .Z(
        n108) );
  OAI21M1P U263 ( .A(n158), .B(n135), .C(n108), .Z(n484) );
  AOI22M1P U264 ( .A(\Queue[2][8] ), .B(n133), .C(n3), .D(\Queue[3][8] ), .Z(
        n109) );
  OAI21M1P U265 ( .A(n160), .B(n135), .C(n109), .Z(n485) );
  AOI22M1P U266 ( .A(\Queue[2][9] ), .B(n133), .C(n3), .D(\Queue[3][9] ), .Z(
        n110) );
  OAI21M1P U267 ( .A(n162), .B(n135), .C(n110), .Z(n486) );
  AOI22M1P U268 ( .A(\Queue[2][10] ), .B(n133), .C(n3), .D(\Queue[3][10] ), 
        .Z(n111) );
  OAI21M1P U269 ( .A(n164), .B(n135), .C(n111), .Z(n487) );
  AOI22M1P U270 ( .A(\Queue[2][11] ), .B(n133), .C(n3), .D(\Queue[3][11] ), 
        .Z(n112) );
  OAI21M1P U271 ( .A(n166), .B(n135), .C(n112), .Z(n488) );
  AOI22M1P U272 ( .A(\Queue[2][12] ), .B(n133), .C(n3), .D(\Queue[3][12] ), 
        .Z(n113) );
  OAI21M1P U273 ( .A(n168), .B(n135), .C(n113), .Z(n489) );
  AOI22M1P U274 ( .A(\Queue[2][13] ), .B(n133), .C(n3), .D(\Queue[3][13] ), 
        .Z(n114) );
  OAI21M1P U275 ( .A(n170), .B(n135), .C(n114), .Z(n490) );
  AOI22M1P U276 ( .A(\Queue[2][14] ), .B(n133), .C(n3), .D(\Queue[3][14] ), 
        .Z(n115) );
  OAI21M1P U277 ( .A(n172), .B(n135), .C(n115), .Z(n491) );
  AOI22M1P U278 ( .A(\Queue[2][15] ), .B(n133), .C(n3), .D(\Queue[3][15] ), 
        .Z(n116) );
  OAI21M1P U279 ( .A(n174), .B(n135), .C(n116), .Z(n492) );
  AOI22M1P U280 ( .A(\Queue[2][16] ), .B(n133), .C(n3), .D(\Queue[3][16] ), 
        .Z(n117) );
  OAI21M1P U281 ( .A(n176), .B(n135), .C(n117), .Z(n493) );
  AOI22M1P U282 ( .A(\Queue[2][17] ), .B(n133), .C(n3), .D(\Queue[3][17] ), 
        .Z(n118) );
  OAI21M1P U283 ( .A(n178), .B(n135), .C(n118), .Z(n494) );
  AOI22M1P U284 ( .A(\Queue[2][18] ), .B(n133), .C(n3), .D(\Queue[3][18] ), 
        .Z(n119) );
  OAI21M1P U285 ( .A(n180), .B(n135), .C(n119), .Z(n495) );
  AOI22M1P U286 ( .A(\Queue[2][19] ), .B(n133), .C(n3), .D(\Queue[3][19] ), 
        .Z(n120) );
  OAI21M1P U287 ( .A(n182), .B(n135), .C(n120), .Z(n496) );
  AOI22M1P U288 ( .A(\Queue[2][20] ), .B(n133), .C(n3), .D(\Queue[3][20] ), 
        .Z(n121) );
  OAI21M1P U289 ( .A(n184), .B(n135), .C(n121), .Z(n497) );
  AOI22M1P U290 ( .A(\Queue[2][21] ), .B(n133), .C(n3), .D(\Queue[3][21] ), 
        .Z(n122) );
  OAI21M1P U291 ( .A(n186), .B(n135), .C(n122), .Z(n498) );
  AOI22M1P U292 ( .A(\Queue[2][22] ), .B(n133), .C(n3), .D(\Queue[3][22] ), 
        .Z(n123) );
  OAI21M1P U293 ( .A(n188), .B(n135), .C(n123), .Z(n499) );
  AOI22M1P U294 ( .A(\Queue[2][23] ), .B(n133), .C(n3), .D(\Queue[3][23] ), 
        .Z(n124) );
  OAI21M1P U295 ( .A(n190), .B(n135), .C(n124), .Z(n500) );
  AOI22M1P U296 ( .A(\Queue[2][24] ), .B(n133), .C(n3), .D(\Queue[3][24] ), 
        .Z(n125) );
  OAI21M1P U297 ( .A(n192), .B(n135), .C(n125), .Z(n501) );
  AOI22M1P U298 ( .A(\Queue[2][25] ), .B(n133), .C(n3), .D(\Queue[3][25] ), 
        .Z(n126) );
  OAI21M1P U299 ( .A(n194), .B(n135), .C(n126), .Z(n502) );
  AOI22M1P U300 ( .A(\Queue[2][26] ), .B(n133), .C(n3), .D(\Queue[3][26] ), 
        .Z(n127) );
  OAI21M1P U301 ( .A(n196), .B(n135), .C(n127), .Z(n503) );
  AOI22M1P U302 ( .A(\Queue[2][27] ), .B(n133), .C(n3), .D(\Queue[3][27] ), 
        .Z(n128) );
  OAI21M1P U303 ( .A(n198), .B(n135), .C(n128), .Z(n504) );
  AOI22M1P U304 ( .A(\Queue[2][28] ), .B(n133), .C(n3), .D(\Queue[3][28] ), 
        .Z(n129) );
  OAI21M1P U305 ( .A(n200), .B(n135), .C(n129), .Z(n505) );
  AOI22M1P U306 ( .A(\Queue[2][29] ), .B(n133), .C(n3), .D(\Queue[3][29] ), 
        .Z(n130) );
  OAI21M1P U307 ( .A(n202), .B(n135), .C(n130), .Z(n506) );
  AOI22M1P U308 ( .A(\Queue[2][30] ), .B(n133), .C(n3), .D(\Queue[3][30] ), 
        .Z(n131) );
  OAI21M1P U309 ( .A(n204), .B(n135), .C(n131), .Z(n507) );
  AOI22M1P U310 ( .A(\Queue[2][31] ), .B(n133), .C(n3), .D(\Queue[3][31] ), 
        .Z(n134) );
  OAI21M1P U311 ( .A(n373), .B(n135), .C(n134), .Z(n508) );
  OA21M1P U312 ( .A(n139), .B(n140), .C(Rst_n), .Z(n136) );
  AOI22M1P U313 ( .A(\Queue[3][0] ), .B(n206), .C(n205), .D(\Queue[4][0] ), 
        .Z(n143) );
  OAI21M1P U314 ( .A(n144), .B(n208), .C(n143), .Z(n509) );
  AOI22M1P U315 ( .A(\Queue[3][1] ), .B(n206), .C(n205), .D(\Queue[4][1] ), 
        .Z(n145) );
  OAI21M1P U316 ( .A(n146), .B(n208), .C(n145), .Z(n510) );
  AOI22M1P U317 ( .A(\Queue[3][2] ), .B(n206), .C(n205), .D(\Queue[4][2] ), 
        .Z(n147) );
  OAI21M1P U318 ( .A(n148), .B(n208), .C(n147), .Z(n511) );
  AOI22M1P U319 ( .A(\Queue[3][3] ), .B(n206), .C(n205), .D(\Queue[4][3] ), 
        .Z(n149) );
  OAI21M1P U320 ( .A(n150), .B(n208), .C(n149), .Z(n512) );
  AOI22M1P U321 ( .A(\Queue[3][4] ), .B(n206), .C(n205), .D(\Queue[4][4] ), 
        .Z(n151) );
  OAI21M1P U322 ( .A(n152), .B(n208), .C(n151), .Z(n513) );
  AOI22M1P U323 ( .A(\Queue[3][5] ), .B(n206), .C(n205), .D(\Queue[4][5] ), 
        .Z(n153) );
  OAI21M1P U324 ( .A(n154), .B(n208), .C(n153), .Z(n514) );
  AOI22M1P U325 ( .A(\Queue[3][6] ), .B(n206), .C(n205), .D(\Queue[4][6] ), 
        .Z(n155) );
  OAI21M1P U326 ( .A(n156), .B(n208), .C(n155), .Z(n515) );
  AOI22M1P U327 ( .A(\Queue[3][7] ), .B(n206), .C(n205), .D(\Queue[4][7] ), 
        .Z(n157) );
  OAI21M1P U328 ( .A(n158), .B(n208), .C(n157), .Z(n516) );
  AOI22M1P U329 ( .A(\Queue[3][8] ), .B(n206), .C(n11), .D(\Queue[4][8] ), .Z(
        n159) );
  OAI21M1P U330 ( .A(n160), .B(n208), .C(n159), .Z(n517) );
  AOI22M1P U331 ( .A(\Queue[3][9] ), .B(n206), .C(n12), .D(\Queue[4][9] ), .Z(
        n161) );
  OAI21M1P U332 ( .A(n162), .B(n208), .C(n161), .Z(n518) );
  AOI22M1P U333 ( .A(\Queue[3][10] ), .B(n206), .C(n11), .D(\Queue[4][10] ), 
        .Z(n163) );
  OAI21M1P U334 ( .A(n164), .B(n208), .C(n163), .Z(n519) );
  AOI22M1P U335 ( .A(\Queue[3][11] ), .B(n206), .C(n11), .D(\Queue[4][11] ), 
        .Z(n165) );
  OAI21M1P U336 ( .A(n166), .B(n208), .C(n165), .Z(n520) );
  AOI22M1P U337 ( .A(\Queue[3][12] ), .B(n206), .C(n11), .D(\Queue[4][12] ), 
        .Z(n167) );
  OAI21M1P U338 ( .A(n168), .B(n208), .C(n167), .Z(n521) );
  AOI22M1P U339 ( .A(\Queue[3][13] ), .B(n206), .C(n11), .D(\Queue[4][13] ), 
        .Z(n169) );
  OAI21M1P U340 ( .A(n170), .B(n208), .C(n169), .Z(n522) );
  AOI22M1P U341 ( .A(\Queue[3][14] ), .B(n206), .C(n11), .D(\Queue[4][14] ), 
        .Z(n171) );
  OAI21M1P U342 ( .A(n172), .B(n208), .C(n171), .Z(n523) );
  AOI22M1P U343 ( .A(\Queue[3][15] ), .B(n206), .C(n11), .D(\Queue[4][15] ), 
        .Z(n173) );
  OAI21M1P U344 ( .A(n174), .B(n208), .C(n173), .Z(n524) );
  AOI22M1P U345 ( .A(\Queue[3][16] ), .B(n206), .C(n11), .D(\Queue[4][16] ), 
        .Z(n175) );
  OAI21M1P U346 ( .A(n176), .B(n208), .C(n175), .Z(n525) );
  AOI22M1P U347 ( .A(\Queue[3][17] ), .B(n206), .C(n11), .D(\Queue[4][17] ), 
        .Z(n177) );
  OAI21M1P U348 ( .A(n178), .B(n208), .C(n177), .Z(n526) );
  AOI22M1P U349 ( .A(\Queue[3][18] ), .B(n206), .C(n11), .D(\Queue[4][18] ), 
        .Z(n179) );
  OAI21M1P U350 ( .A(n180), .B(n208), .C(n179), .Z(n527) );
  AOI22M1P U351 ( .A(\Queue[3][19] ), .B(n206), .C(n11), .D(\Queue[4][19] ), 
        .Z(n181) );
  OAI21M1P U352 ( .A(n182), .B(n208), .C(n181), .Z(n528) );
  AOI22M1P U353 ( .A(\Queue[3][20] ), .B(n206), .C(n12), .D(\Queue[4][20] ), 
        .Z(n183) );
  OAI21M1P U354 ( .A(n184), .B(n208), .C(n183), .Z(n529) );
  AOI22M1P U355 ( .A(\Queue[3][21] ), .B(n206), .C(n12), .D(\Queue[4][21] ), 
        .Z(n185) );
  OAI21M1P U356 ( .A(n186), .B(n208), .C(n185), .Z(n530) );
  AOI22M1P U357 ( .A(\Queue[3][22] ), .B(n206), .C(n12), .D(\Queue[4][22] ), 
        .Z(n187) );
  OAI21M1P U358 ( .A(n188), .B(n208), .C(n187), .Z(n531) );
  AOI22M1P U359 ( .A(\Queue[3][23] ), .B(n206), .C(n12), .D(\Queue[4][23] ), 
        .Z(n189) );
  OAI21M1P U360 ( .A(n190), .B(n208), .C(n189), .Z(n532) );
  AOI22M1P U361 ( .A(\Queue[3][24] ), .B(n206), .C(n12), .D(\Queue[4][24] ), 
        .Z(n191) );
  OAI21M1P U362 ( .A(n192), .B(n208), .C(n191), .Z(n533) );
  AOI22M1P U363 ( .A(\Queue[3][25] ), .B(n206), .C(n12), .D(\Queue[4][25] ), 
        .Z(n193) );
  OAI21M1P U364 ( .A(n194), .B(n208), .C(n193), .Z(n534) );
  AOI22M1P U365 ( .A(\Queue[3][26] ), .B(n206), .C(n12), .D(\Queue[4][26] ), 
        .Z(n195) );
  OAI21M1P U366 ( .A(n196), .B(n208), .C(n195), .Z(n535) );
  AOI22M1P U367 ( .A(\Queue[3][27] ), .B(n206), .C(n12), .D(\Queue[4][27] ), 
        .Z(n197) );
  OAI21M1P U368 ( .A(n198), .B(n208), .C(n197), .Z(n536) );
  AOI22M1P U369 ( .A(\Queue[3][28] ), .B(n206), .C(n12), .D(\Queue[4][28] ), 
        .Z(n199) );
  OAI21M1P U370 ( .A(n200), .B(n208), .C(n199), .Z(n537) );
  AOI22M1P U371 ( .A(\Queue[3][29] ), .B(n206), .C(n12), .D(\Queue[4][29] ), 
        .Z(n201) );
  OAI21M1P U372 ( .A(n202), .B(n208), .C(n201), .Z(n538) );
  AOI22M1P U373 ( .A(\Queue[3][30] ), .B(n206), .C(n11), .D(\Queue[4][30] ), 
        .Z(n203) );
  OAI21M1P U374 ( .A(n204), .B(n208), .C(n203), .Z(n539) );
  AOI22M1P U375 ( .A(\Queue[3][31] ), .B(n206), .C(n12), .D(\Queue[4][31] ), 
        .Z(n207) );
  OAI21M1P U376 ( .A(n373), .B(n208), .C(n207), .Z(n540) );
  N1M1P U377 ( .A(n541), .Z(Empty) );
  AOI22M1P U378 ( .A(n376), .B(n375), .C(n374), .D(Empty), .Z(n542) );
endmodule


module Link_Control_2 ( Clk_r, Rst_n, Tx_Ready, Tx_Error, RxData_Valid, RxData, 
        Packet_From_Core, TxQueue_Write, RxQueue_Read, TxData_Valid, TxData, 
        Error_Ack, Core_Rcv_Ready, Packet_To_Core, RxQueue_Empty, TxQueue_Full
 );
  input [31:0] RxData;
  input [31:0] Packet_From_Core;
  output [31:0] TxData;
  output [31:0] Packet_To_Core;
  input Clk_r, Rst_n, Tx_Ready, Tx_Error, RxData_Valid, TxQueue_Write,
         RxQueue_Read;
  output TxData_Valid, Error_Ack, Core_Rcv_Ready, RxQueue_Empty, TxQueue_Full;
  wire   TxQueue_Read, TxQueue_Empty, RxQueue_Write, RxQueue_Full, N9, N16, n5,
         n6, n7, n8, n9;

  Packet_Queue_6 TxQueue ( .Clk_r(Clk_r), .Rst_n(Rst_n), .Packet_In(
        Packet_From_Core), .Read_Ack(TxQueue_Read), .Write_Ack(TxQueue_Write), 
        .Packet_Out(TxData), .Empty(TxQueue_Empty), .Full(TxQueue_Full) );
  Packet_Queue_5 RxQueue ( .Clk_r(Clk_r), .Rst_n(Rst_n), .Packet_In(RxData), 
        .Read_Ack(RxQueue_Read), .Write_Ack(RxQueue_Write), .Packet_Out(
        Packet_To_Core), .Empty(RxQueue_Empty), .Full(RxQueue_Full) );
  FD2QM1P Core_Rcv_Ready_reg ( .D(N9), .CP(Clk_r), .CD(Rst_n), .Q(
        Core_Rcv_Ready) );
  FD2QM1P TxQueue_Read_reg ( .D(N16), .CP(Clk_r), .CD(Rst_n), .Q(TxQueue_Read)
         );
  FD2QM1P Error_Ack_reg ( .D(Tx_Error), .CP(Clk_r), .CD(Rst_n), .Q(Error_Ack)
         );
  FD4QM1P RxQueue_Write_reg ( .D(n7), .CP(Clk_r), .SD(Rst_n), .Q(n6) );
  FD4QM1P TxData_Valid_reg ( .D(n9), .CP(Clk_r), .SD(Rst_n), .Q(n8) );
  N1M2P U3 ( .A(n6), .Z(RxQueue_Write) );
  NR2M1P U4 ( .A(n8), .B(Tx_Ready), .Z(N16) );
  NR2M1P U5 ( .A(RxData_Valid), .B(RxQueue_Full), .Z(n5) );
  OA21M1P U6 ( .A(Core_Rcv_Ready), .B(n5), .C(n6), .Z(N9) );
  N1M1P U7 ( .A(n8), .Z(TxData_Valid) );
  ND3M1P U8 ( .A(n6), .B(Core_Rcv_Ready), .C(RxData_Valid), .Z(n7) );
  AO21CNM1P U9 ( .A(n8), .B(TxQueue_Empty), .C(Tx_Ready), .Z(n9) );
endmodule


module Packet_Queue_7 ( Clk_r, Rst_n, Packet_In, Read_Ack, Write_Ack, 
        Packet_Out, Empty, Full );
  input [31:0] Packet_In;
  output [31:0] Packet_Out;
  input Clk_r, Rst_n, Read_Ack, Write_Ack;
  output Empty, Full;
  wire   \Queue[4][31] , \Queue[4][30] , \Queue[4][29] , \Queue[4][28] ,
         \Queue[4][27] , \Queue[4][26] , \Queue[4][25] , \Queue[4][24] ,
         \Queue[4][23] , \Queue[4][22] , \Queue[4][21] , \Queue[4][20] ,
         \Queue[4][19] , \Queue[4][18] , \Queue[4][17] , \Queue[4][16] ,
         \Queue[4][15] , \Queue[4][14] , \Queue[4][13] , \Queue[4][12] ,
         \Queue[4][11] , \Queue[4][10] , \Queue[4][9] , \Queue[4][8] ,
         \Queue[4][7] , \Queue[4][6] , \Queue[4][5] , \Queue[4][4] ,
         \Queue[4][3] , \Queue[4][2] , \Queue[4][1] , \Queue[4][0] ,
         \Queue[3][31] , \Queue[3][30] , \Queue[3][29] , \Queue[3][28] ,
         \Queue[3][27] , \Queue[3][26] , \Queue[3][25] , \Queue[3][24] ,
         \Queue[3][23] , \Queue[3][22] , \Queue[3][21] , \Queue[3][20] ,
         \Queue[3][19] , \Queue[3][18] , \Queue[3][17] , \Queue[3][16] ,
         \Queue[3][15] , \Queue[3][14] , \Queue[3][13] , \Queue[3][12] ,
         \Queue[3][11] , \Queue[3][10] , \Queue[3][9] , \Queue[3][8] ,
         \Queue[3][7] , \Queue[3][6] , \Queue[3][5] , \Queue[3][4] ,
         \Queue[3][3] , \Queue[3][2] , \Queue[3][1] , \Queue[3][0] ,
         \Queue[2][31] , \Queue[2][30] , \Queue[2][29] , \Queue[2][28] ,
         \Queue[2][27] , \Queue[2][26] , \Queue[2][25] , \Queue[2][24] ,
         \Queue[2][23] , \Queue[2][22] , \Queue[2][21] , \Queue[2][20] ,
         \Queue[2][19] , \Queue[2][18] , \Queue[2][17] , \Queue[2][16] ,
         \Queue[2][15] , \Queue[2][14] , \Queue[2][13] , \Queue[2][12] ,
         \Queue[2][11] , \Queue[2][10] , \Queue[2][9] , \Queue[2][8] ,
         \Queue[2][7] , \Queue[2][6] , \Queue[2][5] , \Queue[2][4] ,
         \Queue[2][3] , \Queue[2][2] , \Queue[2][1] , \Queue[2][0] ,
         \Queue[1][31] , \Queue[1][30] , \Queue[1][29] , \Queue[1][28] ,
         \Queue[1][27] , \Queue[1][26] , \Queue[1][25] , \Queue[1][24] ,
         \Queue[1][23] , \Queue[1][22] , \Queue[1][21] , \Queue[1][20] ,
         \Queue[1][19] , \Queue[1][18] , \Queue[1][17] , \Queue[1][16] ,
         \Queue[1][15] , \Queue[1][14] , \Queue[1][13] , \Queue[1][12] ,
         \Queue[1][11] , \Queue[1][10] , \Queue[1][9] , \Queue[1][8] ,
         \Queue[1][7] , \Queue[1][6] , \Queue[1][5] , \Queue[1][4] ,
         \Queue[1][3] , \Queue[1][2] , \Queue[1][1] , \Queue[1][0] , n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550;
  wire   [2:0] Count;

  FDN2QM1P \Count_reg[0]  ( .D(n385), .CPN(Clk_r), .CD(Rst_n), .Q(Count[0]) );
  FDN2QM1P \Count_reg[1]  ( .D(n386), .CPN(Clk_r), .CD(Rst_n), .Q(Count[1]) );
  FDN2QM1P \Count_reg[2]  ( .D(n387), .CPN(Clk_r), .CD(Rst_n), .Q(Count[2]) );
  FDN1QM1P \Queue_reg[4][30]  ( .D(n419), .CPN(Clk_r), .Q(\Queue[4][30] ) );
  FDN1QM1P \Queue_reg[3][30]  ( .D(n547), .CPN(Clk_r), .Q(\Queue[3][30] ) );
  FDN1QM1P \Queue_reg[2][30]  ( .D(n515), .CPN(Clk_r), .Q(\Queue[2][30] ) );
  FDN1QM1P \Queue_reg[4][29]  ( .D(n418), .CPN(Clk_r), .Q(\Queue[4][29] ) );
  FDN1QM1P \Queue_reg[3][29]  ( .D(n546), .CPN(Clk_r), .Q(\Queue[3][29] ) );
  FDN1QM1P \Queue_reg[2][29]  ( .D(n514), .CPN(Clk_r), .Q(\Queue[2][29] ) );
  FDN1QM1P \Queue_reg[4][28]  ( .D(n417), .CPN(Clk_r), .Q(\Queue[4][28] ) );
  FDN1QM1P \Queue_reg[3][28]  ( .D(n545), .CPN(Clk_r), .Q(\Queue[3][28] ) );
  FDN1QM1P \Queue_reg[2][28]  ( .D(n513), .CPN(Clk_r), .Q(\Queue[2][28] ) );
  FDN1QM1P \Queue_reg[4][27]  ( .D(n416), .CPN(Clk_r), .Q(\Queue[4][27] ) );
  FDN1QM1P \Queue_reg[3][27]  ( .D(n544), .CPN(Clk_r), .Q(\Queue[3][27] ) );
  FDN1QM1P \Queue_reg[2][27]  ( .D(n512), .CPN(Clk_r), .Q(\Queue[2][27] ) );
  FDN1QM1P \Queue_reg[4][26]  ( .D(n415), .CPN(Clk_r), .Q(\Queue[4][26] ) );
  FDN1QM1P \Queue_reg[3][26]  ( .D(n543), .CPN(Clk_r), .Q(\Queue[3][26] ) );
  FDN1QM1P \Queue_reg[2][26]  ( .D(n511), .CPN(Clk_r), .Q(\Queue[2][26] ) );
  FDN1QM1P \Queue_reg[4][25]  ( .D(n414), .CPN(Clk_r), .Q(\Queue[4][25] ) );
  FDN1QM1P \Queue_reg[3][25]  ( .D(n542), .CPN(Clk_r), .Q(\Queue[3][25] ) );
  FDN1QM1P \Queue_reg[2][25]  ( .D(n510), .CPN(Clk_r), .Q(\Queue[2][25] ) );
  FDN1QM1P \Queue_reg[4][24]  ( .D(n413), .CPN(Clk_r), .Q(\Queue[4][24] ) );
  FDN1QM1P \Queue_reg[3][24]  ( .D(n541), .CPN(Clk_r), .Q(\Queue[3][24] ) );
  FDN1QM1P \Queue_reg[2][24]  ( .D(n509), .CPN(Clk_r), .Q(\Queue[2][24] ) );
  FDN1QM1P \Queue_reg[4][23]  ( .D(n412), .CPN(Clk_r), .Q(\Queue[4][23] ) );
  FDN1QM1P \Queue_reg[3][23]  ( .D(n540), .CPN(Clk_r), .Q(\Queue[3][23] ) );
  FDN1QM1P \Queue_reg[2][23]  ( .D(n508), .CPN(Clk_r), .Q(\Queue[2][23] ) );
  FDN1QM1P \Queue_reg[4][22]  ( .D(n411), .CPN(Clk_r), .Q(\Queue[4][22] ) );
  FDN1QM1P \Queue_reg[3][22]  ( .D(n539), .CPN(Clk_r), .Q(\Queue[3][22] ) );
  FDN1QM1P \Queue_reg[2][22]  ( .D(n507), .CPN(Clk_r), .Q(\Queue[2][22] ) );
  FDN1QM1P \Queue_reg[4][21]  ( .D(n410), .CPN(Clk_r), .Q(\Queue[4][21] ) );
  FDN1QM1P \Queue_reg[3][21]  ( .D(n538), .CPN(Clk_r), .Q(\Queue[3][21] ) );
  FDN1QM1P \Queue_reg[2][21]  ( .D(n506), .CPN(Clk_r), .Q(\Queue[2][21] ) );
  FDN1QM1P \Queue_reg[4][20]  ( .D(n409), .CPN(Clk_r), .Q(\Queue[4][20] ) );
  FDN1QM1P \Queue_reg[3][20]  ( .D(n537), .CPN(Clk_r), .Q(\Queue[3][20] ) );
  FDN1QM1P \Queue_reg[2][20]  ( .D(n505), .CPN(Clk_r), .Q(\Queue[2][20] ) );
  FDN1QM1P \Queue_reg[4][19]  ( .D(n408), .CPN(Clk_r), .Q(\Queue[4][19] ) );
  FDN1QM1P \Queue_reg[3][19]  ( .D(n536), .CPN(Clk_r), .Q(\Queue[3][19] ) );
  FDN1QM1P \Queue_reg[2][19]  ( .D(n504), .CPN(Clk_r), .Q(\Queue[2][19] ) );
  FDN1QM1P \Queue_reg[4][18]  ( .D(n407), .CPN(Clk_r), .Q(\Queue[4][18] ) );
  FDN1QM1P \Queue_reg[3][18]  ( .D(n535), .CPN(Clk_r), .Q(\Queue[3][18] ) );
  FDN1QM1P \Queue_reg[2][18]  ( .D(n503), .CPN(Clk_r), .Q(\Queue[2][18] ) );
  FDN1QM1P \Queue_reg[4][17]  ( .D(n406), .CPN(Clk_r), .Q(\Queue[4][17] ) );
  FDN1QM1P \Queue_reg[3][17]  ( .D(n534), .CPN(Clk_r), .Q(\Queue[3][17] ) );
  FDN1QM1P \Queue_reg[2][17]  ( .D(n502), .CPN(Clk_r), .Q(\Queue[2][17] ) );
  FDN1QM1P \Queue_reg[4][16]  ( .D(n405), .CPN(Clk_r), .Q(\Queue[4][16] ) );
  FDN1QM1P \Queue_reg[3][16]  ( .D(n533), .CPN(Clk_r), .Q(\Queue[3][16] ) );
  FDN1QM1P \Queue_reg[2][16]  ( .D(n501), .CPN(Clk_r), .Q(\Queue[2][16] ) );
  FDN1QM1P \Queue_reg[4][15]  ( .D(n404), .CPN(Clk_r), .Q(\Queue[4][15] ) );
  FDN1QM1P \Queue_reg[3][15]  ( .D(n532), .CPN(Clk_r), .Q(\Queue[3][15] ) );
  FDN1QM1P \Queue_reg[2][15]  ( .D(n500), .CPN(Clk_r), .Q(\Queue[2][15] ) );
  FDN1QM1P \Queue_reg[4][14]  ( .D(n403), .CPN(Clk_r), .Q(\Queue[4][14] ) );
  FDN1QM1P \Queue_reg[3][14]  ( .D(n531), .CPN(Clk_r), .Q(\Queue[3][14] ) );
  FDN1QM1P \Queue_reg[2][14]  ( .D(n499), .CPN(Clk_r), .Q(\Queue[2][14] ) );
  FDN1QM1P \Queue_reg[4][13]  ( .D(n402), .CPN(Clk_r), .Q(\Queue[4][13] ) );
  FDN1QM1P \Queue_reg[3][13]  ( .D(n530), .CPN(Clk_r), .Q(\Queue[3][13] ) );
  FDN1QM1P \Queue_reg[2][13]  ( .D(n498), .CPN(Clk_r), .Q(\Queue[2][13] ) );
  FDN1QM1P \Queue_reg[4][12]  ( .D(n401), .CPN(Clk_r), .Q(\Queue[4][12] ) );
  FDN1QM1P \Queue_reg[3][12]  ( .D(n529), .CPN(Clk_r), .Q(\Queue[3][12] ) );
  FDN1QM1P \Queue_reg[2][12]  ( .D(n497), .CPN(Clk_r), .Q(\Queue[2][12] ) );
  FDN1QM1P \Queue_reg[4][11]  ( .D(n400), .CPN(Clk_r), .Q(\Queue[4][11] ) );
  FDN1QM1P \Queue_reg[3][11]  ( .D(n528), .CPN(Clk_r), .Q(\Queue[3][11] ) );
  FDN1QM1P \Queue_reg[2][11]  ( .D(n496), .CPN(Clk_r), .Q(\Queue[2][11] ) );
  FDN1QM1P \Queue_reg[4][10]  ( .D(n399), .CPN(Clk_r), .Q(\Queue[4][10] ) );
  FDN1QM1P \Queue_reg[3][10]  ( .D(n527), .CPN(Clk_r), .Q(\Queue[3][10] ) );
  FDN1QM1P \Queue_reg[2][10]  ( .D(n495), .CPN(Clk_r), .Q(\Queue[2][10] ) );
  FDN1QM1P \Queue_reg[4][9]  ( .D(n398), .CPN(Clk_r), .Q(\Queue[4][9] ) );
  FDN1QM1P \Queue_reg[3][9]  ( .D(n526), .CPN(Clk_r), .Q(\Queue[3][9] ) );
  FDN1QM1P \Queue_reg[2][9]  ( .D(n494), .CPN(Clk_r), .Q(\Queue[2][9] ) );
  FDN1QM1P \Queue_reg[4][8]  ( .D(n397), .CPN(Clk_r), .Q(\Queue[4][8] ) );
  FDN1QM1P \Queue_reg[3][8]  ( .D(n525), .CPN(Clk_r), .Q(\Queue[3][8] ) );
  FDN1QM1P \Queue_reg[2][8]  ( .D(n493), .CPN(Clk_r), .Q(\Queue[2][8] ) );
  FDN1QM1P \Queue_reg[4][7]  ( .D(n396), .CPN(Clk_r), .Q(\Queue[4][7] ) );
  FDN1QM1P \Queue_reg[3][7]  ( .D(n524), .CPN(Clk_r), .Q(\Queue[3][7] ) );
  FDN1QM1P \Queue_reg[2][7]  ( .D(n492), .CPN(Clk_r), .Q(\Queue[2][7] ) );
  FDN1QM1P \Queue_reg[4][6]  ( .D(n395), .CPN(Clk_r), .Q(\Queue[4][6] ) );
  FDN1QM1P \Queue_reg[3][6]  ( .D(n523), .CPN(Clk_r), .Q(\Queue[3][6] ) );
  FDN1QM1P \Queue_reg[2][6]  ( .D(n491), .CPN(Clk_r), .Q(\Queue[2][6] ) );
  FDN1QM1P \Queue_reg[4][5]  ( .D(n394), .CPN(Clk_r), .Q(\Queue[4][5] ) );
  FDN1QM1P \Queue_reg[3][5]  ( .D(n522), .CPN(Clk_r), .Q(\Queue[3][5] ) );
  FDN1QM1P \Queue_reg[2][5]  ( .D(n490), .CPN(Clk_r), .Q(\Queue[2][5] ) );
  FDN1QM1P \Queue_reg[4][4]  ( .D(n393), .CPN(Clk_r), .Q(\Queue[4][4] ) );
  FDN1QM1P \Queue_reg[3][4]  ( .D(n521), .CPN(Clk_r), .Q(\Queue[3][4] ) );
  FDN1QM1P \Queue_reg[2][4]  ( .D(n489), .CPN(Clk_r), .Q(\Queue[2][4] ) );
  FDN1QM1P \Queue_reg[4][3]  ( .D(n392), .CPN(Clk_r), .Q(\Queue[4][3] ) );
  FDN1QM1P \Queue_reg[3][3]  ( .D(n520), .CPN(Clk_r), .Q(\Queue[3][3] ) );
  FDN1QM1P \Queue_reg[2][3]  ( .D(n488), .CPN(Clk_r), .Q(\Queue[2][3] ) );
  FDN1QM1P \Queue_reg[4][2]  ( .D(n391), .CPN(Clk_r), .Q(\Queue[4][2] ) );
  FDN1QM1P \Queue_reg[3][2]  ( .D(n519), .CPN(Clk_r), .Q(\Queue[3][2] ) );
  FDN1QM1P \Queue_reg[2][2]  ( .D(n487), .CPN(Clk_r), .Q(\Queue[2][2] ) );
  FDN1QM1P \Queue_reg[4][1]  ( .D(n390), .CPN(Clk_r), .Q(\Queue[4][1] ) );
  FDN1QM1P \Queue_reg[3][1]  ( .D(n518), .CPN(Clk_r), .Q(\Queue[3][1] ) );
  FDN1QM1P \Queue_reg[2][1]  ( .D(n486), .CPN(Clk_r), .Q(\Queue[2][1] ) );
  FDN1QM1P \Queue_reg[4][0]  ( .D(n389), .CPN(Clk_r), .Q(\Queue[4][0] ) );
  FDN1QM1P \Queue_reg[3][0]  ( .D(n517), .CPN(Clk_r), .Q(\Queue[3][0] ) );
  FDN1QM1P \Queue_reg[4][31]  ( .D(n388), .CPN(Clk_r), .Q(\Queue[4][31] ) );
  FDN1QM1P \Queue_reg[3][31]  ( .D(n548), .CPN(Clk_r), .Q(\Queue[3][31] ) );
  FDN1QM1P \Queue_reg[2][31]  ( .D(n516), .CPN(Clk_r), .Q(\Queue[2][31] ) );
  FDN2QM1P Full_reg ( .D(n420), .CPN(Clk_r), .CD(Rst_n), .Q(Full) );
  FDN1QM1P \Queue_reg[1][31]  ( .D(n452), .CPN(Clk_r), .Q(\Queue[1][31] ) );
  FDN1QM1P \Queue_reg[0][31]  ( .D(n484), .CPN(Clk_r), .Q(Packet_Out[31]) );
  FDN1QM1P \Queue_reg[1][30]  ( .D(n451), .CPN(Clk_r), .Q(\Queue[1][30] ) );
  FDN1QM1P \Queue_reg[0][30]  ( .D(n483), .CPN(Clk_r), .Q(Packet_Out[30]) );
  FDN1QM1P \Queue_reg[1][29]  ( .D(n450), .CPN(Clk_r), .Q(\Queue[1][29] ) );
  FDN1QM1P \Queue_reg[0][29]  ( .D(n482), .CPN(Clk_r), .Q(Packet_Out[29]) );
  FDN1QM1P \Queue_reg[1][28]  ( .D(n449), .CPN(Clk_r), .Q(\Queue[1][28] ) );
  FDN1QM1P \Queue_reg[0][28]  ( .D(n481), .CPN(Clk_r), .Q(Packet_Out[28]) );
  FDN1QM1P \Queue_reg[1][27]  ( .D(n448), .CPN(Clk_r), .Q(\Queue[1][27] ) );
  FDN1QM1P \Queue_reg[0][27]  ( .D(n480), .CPN(Clk_r), .Q(Packet_Out[27]) );
  FDN1QM1P \Queue_reg[1][26]  ( .D(n447), .CPN(Clk_r), .Q(\Queue[1][26] ) );
  FDN1QM1P \Queue_reg[0][26]  ( .D(n479), .CPN(Clk_r), .Q(Packet_Out[26]) );
  FDN1QM1P \Queue_reg[1][25]  ( .D(n446), .CPN(Clk_r), .Q(\Queue[1][25] ) );
  FDN1QM1P \Queue_reg[0][25]  ( .D(n478), .CPN(Clk_r), .Q(Packet_Out[25]) );
  FDN1QM1P \Queue_reg[1][24]  ( .D(n445), .CPN(Clk_r), .Q(\Queue[1][24] ) );
  FDN1QM1P \Queue_reg[0][24]  ( .D(n477), .CPN(Clk_r), .Q(Packet_Out[24]) );
  FDN1QM1P \Queue_reg[1][23]  ( .D(n444), .CPN(Clk_r), .Q(\Queue[1][23] ) );
  FDN1QM1P \Queue_reg[0][23]  ( .D(n476), .CPN(Clk_r), .Q(Packet_Out[23]) );
  FDN1QM1P \Queue_reg[1][22]  ( .D(n443), .CPN(Clk_r), .Q(\Queue[1][22] ) );
  FDN1QM1P \Queue_reg[0][22]  ( .D(n475), .CPN(Clk_r), .Q(Packet_Out[22]) );
  FDN1QM1P \Queue_reg[1][21]  ( .D(n442), .CPN(Clk_r), .Q(\Queue[1][21] ) );
  FDN1QM1P \Queue_reg[0][21]  ( .D(n474), .CPN(Clk_r), .Q(Packet_Out[21]) );
  FDN1QM1P \Queue_reg[1][20]  ( .D(n441), .CPN(Clk_r), .Q(\Queue[1][20] ) );
  FDN1QM1P \Queue_reg[0][20]  ( .D(n473), .CPN(Clk_r), .Q(Packet_Out[20]) );
  FDN1QM1P \Queue_reg[1][19]  ( .D(n440), .CPN(Clk_r), .Q(\Queue[1][19] ) );
  FDN1QM1P \Queue_reg[0][19]  ( .D(n472), .CPN(Clk_r), .Q(Packet_Out[19]) );
  FDN1QM1P \Queue_reg[1][18]  ( .D(n439), .CPN(Clk_r), .Q(\Queue[1][18] ) );
  FDN1QM1P \Queue_reg[0][18]  ( .D(n471), .CPN(Clk_r), .Q(Packet_Out[18]) );
  FDN1QM1P \Queue_reg[1][17]  ( .D(n438), .CPN(Clk_r), .Q(\Queue[1][17] ) );
  FDN1QM1P \Queue_reg[0][17]  ( .D(n470), .CPN(Clk_r), .Q(Packet_Out[17]) );
  FDN1QM1P \Queue_reg[1][16]  ( .D(n437), .CPN(Clk_r), .Q(\Queue[1][16] ) );
  FDN1QM1P \Queue_reg[0][16]  ( .D(n469), .CPN(Clk_r), .Q(Packet_Out[16]) );
  FDN1QM1P \Queue_reg[1][15]  ( .D(n436), .CPN(Clk_r), .Q(\Queue[1][15] ) );
  FDN1QM1P \Queue_reg[0][15]  ( .D(n468), .CPN(Clk_r), .Q(Packet_Out[15]) );
  FDN1QM1P \Queue_reg[1][14]  ( .D(n435), .CPN(Clk_r), .Q(\Queue[1][14] ) );
  FDN1QM1P \Queue_reg[0][14]  ( .D(n467), .CPN(Clk_r), .Q(Packet_Out[14]) );
  FDN1QM1P \Queue_reg[1][13]  ( .D(n434), .CPN(Clk_r), .Q(\Queue[1][13] ) );
  FDN1QM1P \Queue_reg[0][13]  ( .D(n466), .CPN(Clk_r), .Q(Packet_Out[13]) );
  FDN1QM1P \Queue_reg[1][12]  ( .D(n433), .CPN(Clk_r), .Q(\Queue[1][12] ) );
  FDN1QM1P \Queue_reg[0][12]  ( .D(n465), .CPN(Clk_r), .Q(Packet_Out[12]) );
  FDN1QM1P \Queue_reg[1][11]  ( .D(n432), .CPN(Clk_r), .Q(\Queue[1][11] ) );
  FDN1QM1P \Queue_reg[0][11]  ( .D(n464), .CPN(Clk_r), .Q(Packet_Out[11]) );
  FDN1QM1P \Queue_reg[1][10]  ( .D(n431), .CPN(Clk_r), .Q(\Queue[1][10] ) );
  FDN1QM1P \Queue_reg[0][10]  ( .D(n463), .CPN(Clk_r), .Q(Packet_Out[10]) );
  FDN1QM1P \Queue_reg[1][9]  ( .D(n430), .CPN(Clk_r), .Q(\Queue[1][9] ) );
  FDN1QM1P \Queue_reg[0][9]  ( .D(n462), .CPN(Clk_r), .Q(Packet_Out[9]) );
  FDN1QM1P \Queue_reg[1][8]  ( .D(n429), .CPN(Clk_r), .Q(\Queue[1][8] ) );
  FDN1QM1P \Queue_reg[0][8]  ( .D(n461), .CPN(Clk_r), .Q(Packet_Out[8]) );
  FDN1QM1P \Queue_reg[1][7]  ( .D(n428), .CPN(Clk_r), .Q(\Queue[1][7] ) );
  FDN1QM1P \Queue_reg[0][7]  ( .D(n460), .CPN(Clk_r), .Q(Packet_Out[7]) );
  FDN1QM1P \Queue_reg[1][6]  ( .D(n427), .CPN(Clk_r), .Q(\Queue[1][6] ) );
  FDN1QM1P \Queue_reg[0][6]  ( .D(n459), .CPN(Clk_r), .Q(Packet_Out[6]) );
  FDN1QM1P \Queue_reg[1][5]  ( .D(n426), .CPN(Clk_r), .Q(\Queue[1][5] ) );
  FDN1QM1P \Queue_reg[0][5]  ( .D(n458), .CPN(Clk_r), .Q(Packet_Out[5]) );
  FDN1QM1P \Queue_reg[1][4]  ( .D(n425), .CPN(Clk_r), .Q(\Queue[1][4] ) );
  FDN1QM1P \Queue_reg[0][4]  ( .D(n457), .CPN(Clk_r), .Q(Packet_Out[4]) );
  FDN1QM1P \Queue_reg[1][3]  ( .D(n424), .CPN(Clk_r), .Q(\Queue[1][3] ) );
  FDN1QM1P \Queue_reg[0][3]  ( .D(n456), .CPN(Clk_r), .Q(Packet_Out[3]) );
  FDN1QM1P \Queue_reg[1][2]  ( .D(n423), .CPN(Clk_r), .Q(\Queue[1][2] ) );
  FDN1QM1P \Queue_reg[0][2]  ( .D(n455), .CPN(Clk_r), .Q(Packet_Out[2]) );
  FDN1QM1P \Queue_reg[1][1]  ( .D(n422), .CPN(Clk_r), .Q(\Queue[1][1] ) );
  FDN1QM1P \Queue_reg[0][1]  ( .D(n454), .CPN(Clk_r), .Q(Packet_Out[1]) );
  FDN1QM1P \Queue_reg[1][0]  ( .D(n421), .CPN(Clk_r), .Q(\Queue[1][0] ) );
  FDN1QM1P \Queue_reg[0][0]  ( .D(n453), .CPN(Clk_r), .Q(Packet_Out[0]) );
  FDN2QM1P Empty_reg ( .D(n550), .CPN(Clk_r), .CD(Rst_n), .Q(n549) );
  FDN1QM1P \Queue_reg[2][0]  ( .D(n485), .CPN(Clk_r), .Q(\Queue[2][0] ) );
  NR3M1P U3 ( .A(Count[0]), .B(Count[2]), .C(n63), .Z(n140) );
  BUFM1P U4 ( .A(n100), .Z(n48) );
  N1M2P U5 ( .A(n103), .Z(n135) );
  N1M8P U6 ( .A(n3), .Z(n4) );
  N1M3P U7 ( .A(n138), .Z(n3) );
  OAI211M1P U8 ( .A(n384), .B(n146), .C(Write_Ack), .D(n103), .Z(n138) );
  BUFM1P U9 ( .A(n97), .Z(n44) );
  BUFM2P U10 ( .A(n100), .Z(n47) );
  BUFM2P U11 ( .A(n143), .Z(n50) );
  BUFM1P U12 ( .A(n143), .Z(n49) );
  ND2M2P U13 ( .A(n11), .B(n10), .Z(n52) );
  NR3M1P U14 ( .A(n64), .B(Count[2]), .C(Count[1]), .Z(n384) );
  N1M1P U15 ( .A(Read_Ack), .Z(n146) );
  OAI211M1P U16 ( .A(n149), .B(n148), .C(Rst_n), .D(n147), .Z(n378) );
  NR3M1P U17 ( .A(Count[2]), .B(n64), .C(n63), .Z(n149) );
  BUFM6P U18 ( .A(n144), .Z(n51) );
  N1M4P U19 ( .A(n59), .Z(n148) );
  BUFM8P U20 ( .A(n378), .Z(n53) );
  BUFM1P U21 ( .A(n98), .Z(n46) );
  BUFM1P U22 ( .A(n98), .Z(n45) );
  ND2BNM2P U23 ( .B(n7), .A(n8), .Z(n380) );
  N1M1P U24 ( .A(n61), .Z(n6) );
  N1M2P U25 ( .A(n6), .Z(n5) );
  N1M2P U26 ( .A(n6), .Z(n41) );
  NR2M3P U27 ( .A(n139), .B(Read_Ack), .Z(n59) );
  NR3M1P U28 ( .A(Count[0]), .B(Count[1]), .C(n60), .Z(n151) );
  N1M1P U29 ( .A(n151), .Z(n62) );
  N1M1P U30 ( .A(Count[2]), .Z(n60) );
  N1M1P U31 ( .A(Count[1]), .Z(n63) );
  N1M1P U32 ( .A(Count[0]), .Z(n64) );
  NR2FM2P U33 ( .A(n102), .B(n62), .Z(n61) );
  AOI21M6P U34 ( .A(Write_Ack), .B(n384), .C(n150), .Z(n136) );
  OAI21M1P U35 ( .A(n102), .B(n101), .C(n150), .Z(n103) );
  N1M4P U36 ( .A(Write_Ack), .Z(n139) );
  OAI21M2P U37 ( .A(Write_Ack), .B(Read_Ack), .C(n65), .Z(n97) );
  N1M1P U38 ( .A(Packet_In[1]), .Z(n154) );
  N1M1P U39 ( .A(Packet_In[2]), .Z(n156) );
  N1M1P U40 ( .A(Packet_In[5]), .Z(n162) );
  N1M1P U41 ( .A(Packet_In[4]), .Z(n160) );
  N1M1P U42 ( .A(Packet_In[3]), .Z(n158) );
  N1M1P U43 ( .A(Packet_In[7]), .Z(n166) );
  N1M1P U44 ( .A(Packet_In[6]), .Z(n164) );
  N1M1P U45 ( .A(Packet_In[8]), .Z(n168) );
  N1M1P U46 ( .A(Packet_In[19]), .Z(n190) );
  N1M1P U47 ( .A(Packet_In[10]), .Z(n172) );
  N1M1P U48 ( .A(Packet_In[11]), .Z(n174) );
  N1M1P U49 ( .A(Packet_In[15]), .Z(n182) );
  N1M1P U50 ( .A(Packet_In[9]), .Z(n170) );
  N1M1P U51 ( .A(Packet_In[20]), .Z(n192) );
  N1M1P U52 ( .A(Packet_In[17]), .Z(n186) );
  N1M1P U53 ( .A(Packet_In[13]), .Z(n178) );
  N1M1P U54 ( .A(Packet_In[0]), .Z(n152) );
  N1M1P U55 ( .A(Packet_In[23]), .Z(n198) );
  N1M1P U56 ( .A(Packet_In[21]), .Z(n194) );
  N1M1P U57 ( .A(Packet_In[24]), .Z(n200) );
  N1M1P U58 ( .A(Packet_In[30]), .Z(n376) );
  N1M1P U59 ( .A(Packet_In[22]), .Z(n196) );
  N1M1P U60 ( .A(Packet_In[29]), .Z(n374) );
  N1M1P U61 ( .A(Packet_In[31]), .Z(n381) );
  N1M1P U62 ( .A(Packet_In[26]), .Z(n204) );
  N1M1P U63 ( .A(Packet_In[18]), .Z(n188) );
  N1M1P U64 ( .A(Packet_In[27]), .Z(n206) );
  N1M1P U65 ( .A(Packet_In[12]), .Z(n176) );
  N1M1P U66 ( .A(Packet_In[25]), .Z(n202) );
  N1M1P U67 ( .A(Packet_In[14]), .Z(n180) );
  N1M1P U68 ( .A(Packet_In[28]), .Z(n208) );
  ND2M2P U69 ( .A(Read_Ack), .B(Rst_n), .Z(n150) );
  N1M1P U70 ( .A(Packet_In[16]), .Z(n184) );
  AOI21M6P U71 ( .A(Write_Ack), .B(n151), .C(n150), .Z(n377) );
  ND2M2P U72 ( .A(n59), .B(Rst_n), .Z(n102) );
  BUFM2P U73 ( .A(n97), .Z(n43) );
  BUFM2P U74 ( .A(n97), .Z(n42) );
  OAI211M1P U75 ( .A(n140), .B(n146), .C(Write_Ack), .D(n65), .Z(n100) );
  ND2BNM1P U76 ( .B(n149), .A(n59), .Z(n8) );
  OAI21M1P U77 ( .A(n152), .B(n47), .C(n66), .Z(n421) );
  AOI22M1P U78 ( .A(\Queue[2][0] ), .B(n45), .C(\Queue[1][0] ), .D(n44), .Z(
        n66) );
  OAI211M1P U79 ( .A(n151), .B(n146), .C(Rst_n), .D(Write_Ack), .Z(n7) );
  OAI211M1P U80 ( .A(n140), .B(n148), .C(Rst_n), .D(n147), .Z(n144) );
  AOI22M1P U81 ( .A(\Queue[3][0] ), .B(n53), .C(n377), .D(\Queue[4][0] ), .Z(
        n9) );
  OAI21M1P U82 ( .A(n152), .B(n380), .C(n9), .Z(n517) );
  OA21M1P U83 ( .A(n149), .B(n146), .C(Write_Ack), .Z(n10) );
  OAI21M1P U84 ( .A(n182), .B(n52), .C(n12), .Z(n500) );
  OAI21M1P U85 ( .A(n180), .B(n52), .C(n14), .Z(n499) );
  OAI21M1P U86 ( .A(n178), .B(n52), .C(n18), .Z(n498) );
  OAI21M1P U87 ( .A(n176), .B(n52), .C(n21), .Z(n497) );
  OAI21M1P U88 ( .A(n174), .B(n52), .C(n26), .Z(n496) );
  OAI21M1P U89 ( .A(n172), .B(n52), .C(n29), .Z(n495) );
  OAI21M1P U90 ( .A(n190), .B(n52), .C(n31), .Z(n504) );
  OAI21M1P U91 ( .A(n188), .B(n52), .C(n32), .Z(n503) );
  OAI21M1P U92 ( .A(n186), .B(n52), .C(n34), .Z(n502) );
  OAI21M1P U93 ( .A(n184), .B(n52), .C(n35), .Z(n501) );
  OAI21M1P U94 ( .A(n166), .B(n52), .C(n15), .Z(n492) );
  OAI21M1P U95 ( .A(n164), .B(n52), .C(n22), .Z(n491) );
  OAI21M1P U96 ( .A(n158), .B(n52), .C(n23), .Z(n488) );
  OAI21M1P U97 ( .A(n162), .B(n52), .C(n30), .Z(n490) );
  OAI21M1P U98 ( .A(n170), .B(n52), .C(n33), .Z(n494) );
  OAI21M1P U99 ( .A(n168), .B(n52), .C(n36), .Z(n493) );
  OAI21M1P U100 ( .A(n160), .B(n52), .C(n37), .Z(n489) );
  OAI21M1P U101 ( .A(n156), .B(n52), .C(n38), .Z(n487) );
  OAI21M1P U102 ( .A(n154), .B(n52), .C(n40), .Z(n486) );
  OAI21M1P U103 ( .A(n152), .B(n52), .C(n141), .Z(n485) );
  OAI21M1P U104 ( .A(n208), .B(n52), .C(n13), .Z(n513) );
  OAI21M1P U105 ( .A(n206), .B(n52), .C(n16), .Z(n512) );
  OAI21M1P U106 ( .A(n204), .B(n52), .C(n17), .Z(n511) );
  OAI21M1P U107 ( .A(n202), .B(n52), .C(n19), .Z(n510) );
  OAI21M1P U108 ( .A(n200), .B(n52), .C(n20), .Z(n509) );
  OAI21M1P U109 ( .A(n198), .B(n52), .C(n24), .Z(n508) );
  OAI21M1P U110 ( .A(n196), .B(n52), .C(n25), .Z(n507) );
  OAI21M1P U111 ( .A(n194), .B(n52), .C(n27), .Z(n506) );
  OAI21M1P U112 ( .A(n192), .B(n52), .C(n28), .Z(n505) );
  OAI21M1P U113 ( .A(n374), .B(n52), .C(n39), .Z(n514) );
  OA21M1P U114 ( .A(n148), .B(n140), .C(Rst_n), .Z(n11) );
  AOI22M1P U115 ( .A(\Queue[2][15] ), .B(n51), .C(n50), .D(\Queue[3][15] ), 
        .Z(n12) );
  AOI22M1P U116 ( .A(\Queue[2][28] ), .B(n51), .C(n49), .D(\Queue[3][28] ), 
        .Z(n13) );
  AOI22M1P U117 ( .A(\Queue[2][14] ), .B(n51), .C(n50), .D(\Queue[3][14] ), 
        .Z(n14) );
  AOI22M1P U118 ( .A(\Queue[2][7] ), .B(n51), .C(n50), .D(\Queue[3][7] ), .Z(
        n15) );
  AOI22M1P U119 ( .A(\Queue[2][27] ), .B(n51), .C(n49), .D(\Queue[3][27] ), 
        .Z(n16) );
  AOI22M1P U120 ( .A(\Queue[2][26] ), .B(n51), .C(n49), .D(\Queue[3][26] ), 
        .Z(n17) );
  AOI22M1P U121 ( .A(\Queue[2][13] ), .B(n51), .C(n50), .D(\Queue[3][13] ), 
        .Z(n18) );
  AOI22M1P U122 ( .A(\Queue[2][25] ), .B(n51), .C(n49), .D(\Queue[3][25] ), 
        .Z(n19) );
  AOI22M1P U123 ( .A(\Queue[2][24] ), .B(n51), .C(n49), .D(\Queue[3][24] ), 
        .Z(n20) );
  AOI22M1P U124 ( .A(\Queue[2][12] ), .B(n51), .C(n50), .D(\Queue[3][12] ), 
        .Z(n21) );
  AOI22M1P U125 ( .A(\Queue[2][6] ), .B(n51), .C(n50), .D(\Queue[3][6] ), .Z(
        n22) );
  AOI22M1P U126 ( .A(\Queue[2][3] ), .B(n51), .C(n50), .D(\Queue[3][3] ), .Z(
        n23) );
  AOI22M1P U127 ( .A(\Queue[2][23] ), .B(n144), .C(n49), .D(\Queue[3][23] ), 
        .Z(n24) );
  AOI22M1P U128 ( .A(\Queue[2][22] ), .B(n144), .C(n49), .D(\Queue[3][22] ), 
        .Z(n25) );
  AOI22M1P U129 ( .A(\Queue[2][11] ), .B(n51), .C(n50), .D(\Queue[3][11] ), 
        .Z(n26) );
  AOI22M1P U130 ( .A(\Queue[2][21] ), .B(n51), .C(n50), .D(\Queue[3][21] ), 
        .Z(n27) );
  AOI22M1P U131 ( .A(\Queue[2][20] ), .B(n51), .C(n50), .D(\Queue[3][20] ), 
        .Z(n28) );
  AOI22M1P U132 ( .A(\Queue[2][10] ), .B(n51), .C(n50), .D(\Queue[3][10] ), 
        .Z(n29) );
  AOI22M1P U133 ( .A(\Queue[2][5] ), .B(n51), .C(n50), .D(\Queue[3][5] ), .Z(
        n30) );
  AOI22M1P U134 ( .A(\Queue[2][19] ), .B(n51), .C(n50), .D(\Queue[3][19] ), 
        .Z(n31) );
  AOI22M1P U135 ( .A(\Queue[2][18] ), .B(n51), .C(n50), .D(\Queue[3][18] ), 
        .Z(n32) );
  AOI22M1P U136 ( .A(\Queue[2][9] ), .B(n51), .C(n50), .D(\Queue[3][9] ), .Z(
        n33) );
  AOI22M1P U137 ( .A(\Queue[2][17] ), .B(n51), .C(n50), .D(\Queue[3][17] ), 
        .Z(n34) );
  AOI22M1P U138 ( .A(\Queue[2][16] ), .B(n51), .C(n50), .D(\Queue[3][16] ), 
        .Z(n35) );
  AOI22M1P U139 ( .A(\Queue[2][8] ), .B(n51), .C(n50), .D(\Queue[3][8] ), .Z(
        n36) );
  AOI22M1P U140 ( .A(\Queue[2][4] ), .B(n51), .C(n50), .D(\Queue[3][4] ), .Z(
        n37) );
  AOI22M1P U141 ( .A(\Queue[2][2] ), .B(n51), .C(n50), .D(\Queue[3][2] ), .Z(
        n38) );
  AOI22M1P U142 ( .A(\Queue[2][29] ), .B(n144), .C(n49), .D(\Queue[3][29] ), 
        .Z(n39) );
  AOI22M1P U143 ( .A(\Queue[2][1] ), .B(n51), .C(n49), .D(\Queue[3][1] ), .Z(
        n40) );
  NR2M1P U144 ( .A(n146), .B(Write_Ack), .Z(n383) );
  NR2M1P U145 ( .A(n59), .B(n383), .Z(n382) );
  AOI22CDNM1P U146 ( .A(n382), .B(n64), .C(n382), .D(n64), .Z(n385) );
  N1M1P U147 ( .A(n383), .Z(n58) );
  AOI22M1P U148 ( .A(Count[0]), .B(n148), .C(n58), .D(n64), .Z(n55) );
  AOI22CDNM1P U149 ( .A(Count[1]), .B(n55), .C(n55), .D(Count[1]), .Z(n386) );
  ND3M1P U150 ( .A(n64), .B(n60), .C(n63), .Z(n101) );
  ND2M1P U151 ( .A(Count[1]), .B(Read_Ack), .Z(n54) );
  OAI211M1P U152 ( .A(Count[1]), .B(n148), .C(n55), .D(n54), .Z(n56) );
  AOI22M1P U153 ( .A(n59), .B(n149), .C(Count[2]), .D(n56), .Z(n57) );
  OAI21M1P U154 ( .A(n101), .B(n58), .C(n57), .Z(n387) );
  AOI22CDNM1P U155 ( .A(n5), .B(n381), .C(\Queue[4][31] ), .D(n61), .Z(n388)
         );
  AOI22CDNM1P U156 ( .A(n5), .B(n152), .C(\Queue[4][0] ), .D(n41), .Z(n389) );
  AOI22CDNM1P U157 ( .A(n5), .B(n154), .C(\Queue[4][1] ), .D(n41), .Z(n390) );
  AOI22CDNM1P U158 ( .A(n5), .B(n156), .C(\Queue[4][2] ), .D(n41), .Z(n391) );
  AOI22CDNM1P U159 ( .A(n5), .B(n158), .C(\Queue[4][3] ), .D(n41), .Z(n392) );
  AOI22CDNM1P U160 ( .A(n5), .B(n160), .C(\Queue[4][4] ), .D(n41), .Z(n393) );
  AOI22CDNM1P U161 ( .A(n5), .B(n162), .C(\Queue[4][5] ), .D(n41), .Z(n394) );
  AOI22CDNM1P U162 ( .A(n5), .B(n164), .C(\Queue[4][6] ), .D(n5), .Z(n395) );
  AOI22CDNM1P U163 ( .A(n5), .B(n166), .C(\Queue[4][7] ), .D(n5), .Z(n396) );
  AOI22CDNM1P U164 ( .A(n5), .B(n168), .C(\Queue[4][8] ), .D(n41), .Z(n397) );
  AOI22CDNM1P U165 ( .A(n5), .B(n170), .C(\Queue[4][9] ), .D(n5), .Z(n398) );
  AOI22CDNM1P U166 ( .A(n5), .B(n172), .C(\Queue[4][10] ), .D(n5), .Z(n399) );
  AOI22CDNM1P U167 ( .A(n5), .B(n174), .C(\Queue[4][11] ), .D(n5), .Z(n400) );
  AOI22CDNM1P U168 ( .A(n5), .B(n176), .C(\Queue[4][12] ), .D(n5), .Z(n401) );
  AOI22CDNM1P U169 ( .A(n5), .B(n178), .C(\Queue[4][13] ), .D(n5), .Z(n402) );
  AOI22CDNM1P U170 ( .A(n5), .B(n180), .C(\Queue[4][14] ), .D(n41), .Z(n403)
         );
  AOI22CDNM1P U171 ( .A(n5), .B(n182), .C(\Queue[4][15] ), .D(n5), .Z(n404) );
  AOI22CDNM1P U172 ( .A(n5), .B(n184), .C(\Queue[4][16] ), .D(n5), .Z(n405) );
  AOI22CDNM1P U173 ( .A(n5), .B(n186), .C(\Queue[4][17] ), .D(n41), .Z(n406)
         );
  AOI22CDNM1P U174 ( .A(n5), .B(n188), .C(\Queue[4][18] ), .D(n41), .Z(n407)
         );
  AOI22CDNM1P U175 ( .A(n5), .B(n190), .C(\Queue[4][19] ), .D(n41), .Z(n408)
         );
  AOI22CDNM1P U176 ( .A(n41), .B(n192), .C(\Queue[4][20] ), .D(n41), .Z(n409)
         );
  AOI22CDNM1P U177 ( .A(n41), .B(n194), .C(\Queue[4][21] ), .D(n41), .Z(n410)
         );
  AOI22CDNM1P U178 ( .A(n41), .B(n196), .C(\Queue[4][22] ), .D(n41), .Z(n411)
         );
  AOI22CDNM1P U179 ( .A(n41), .B(n198), .C(\Queue[4][23] ), .D(n41), .Z(n412)
         );
  AOI22CDNM1P U180 ( .A(n41), .B(n200), .C(\Queue[4][24] ), .D(n41), .Z(n413)
         );
  AOI22CDNM1P U181 ( .A(n41), .B(n202), .C(\Queue[4][25] ), .D(n41), .Z(n414)
         );
  AOI22CDNM1P U182 ( .A(n41), .B(n204), .C(\Queue[4][26] ), .D(n41), .Z(n415)
         );
  AOI22CDNM1P U183 ( .A(n41), .B(n206), .C(\Queue[4][27] ), .D(n41), .Z(n416)
         );
  AOI22CDNM1P U184 ( .A(n41), .B(n208), .C(\Queue[4][28] ), .D(n41), .Z(n417)
         );
  AOI22CDNM1P U185 ( .A(n41), .B(n374), .C(\Queue[4][29] ), .D(n41), .Z(n418)
         );
  AOI22CDNM1P U186 ( .A(n5), .B(n376), .C(\Queue[4][30] ), .D(n41), .Z(n419)
         );
  OAI22CDNM1P U187 ( .A(n148), .B(n62), .C(n382), .D(Full), .Z(n420) );
  OA21M1P U188 ( .A(n148), .B(n384), .C(Rst_n), .Z(n65) );
  AOI21M1P U189 ( .A(Write_Ack), .B(n140), .C(n150), .Z(n98) );
  AOI22M1P U190 ( .A(n46), .B(\Queue[2][1] ), .C(\Queue[1][1] ), .D(n97), .Z(
        n67) );
  OAI21M1P U191 ( .A(n48), .B(n154), .C(n67), .Z(n422) );
  AOI22M1P U192 ( .A(n46), .B(\Queue[2][2] ), .C(\Queue[1][2] ), .D(n97), .Z(
        n68) );
  OAI21M1P U193 ( .A(n48), .B(n156), .C(n68), .Z(n423) );
  AOI22M1P U194 ( .A(n46), .B(\Queue[2][3] ), .C(\Queue[1][3] ), .D(n97), .Z(
        n69) );
  OAI21M1P U195 ( .A(n48), .B(n158), .C(n69), .Z(n424) );
  AOI22M1P U196 ( .A(n46), .B(\Queue[2][4] ), .C(\Queue[1][4] ), .D(n97), .Z(
        n70) );
  OAI21M1P U197 ( .A(n48), .B(n160), .C(n70), .Z(n425) );
  AOI22M1P U198 ( .A(n46), .B(\Queue[2][5] ), .C(\Queue[1][5] ), .D(n42), .Z(
        n71) );
  OAI21M1P U199 ( .A(n48), .B(n162), .C(n71), .Z(n426) );
  AOI22M1P U200 ( .A(n46), .B(\Queue[2][6] ), .C(\Queue[1][6] ), .D(n43), .Z(
        n72) );
  OAI21M1P U201 ( .A(n48), .B(n164), .C(n72), .Z(n427) );
  AOI22M1P U202 ( .A(n46), .B(\Queue[2][7] ), .C(\Queue[1][7] ), .D(n42), .Z(
        n73) );
  OAI21M1P U203 ( .A(n48), .B(n166), .C(n73), .Z(n428) );
  AOI22M1P U204 ( .A(n46), .B(\Queue[2][8] ), .C(\Queue[1][8] ), .D(n43), .Z(
        n74) );
  OAI21M1P U205 ( .A(n48), .B(n168), .C(n74), .Z(n429) );
  AOI22M1P U206 ( .A(n46), .B(\Queue[2][9] ), .C(\Queue[1][9] ), .D(n42), .Z(
        n75) );
  OAI21M1P U207 ( .A(n48), .B(n170), .C(n75), .Z(n430) );
  AOI22M1P U208 ( .A(n46), .B(\Queue[2][10] ), .C(\Queue[1][10] ), .D(n42), 
        .Z(n76) );
  OAI21M1P U209 ( .A(n48), .B(n172), .C(n76), .Z(n431) );
  AOI22M1P U210 ( .A(n46), .B(\Queue[2][11] ), .C(\Queue[1][11] ), .D(n42), 
        .Z(n77) );
  OAI21M1P U211 ( .A(n48), .B(n174), .C(n77), .Z(n432) );
  AOI22M1P U212 ( .A(n45), .B(\Queue[2][12] ), .C(\Queue[1][12] ), .D(n42), 
        .Z(n78) );
  OAI21M1P U213 ( .A(n47), .B(n176), .C(n78), .Z(n433) );
  AOI22M1P U214 ( .A(n46), .B(\Queue[2][13] ), .C(\Queue[1][13] ), .D(n42), 
        .Z(n79) );
  OAI21M1P U215 ( .A(n47), .B(n178), .C(n79), .Z(n434) );
  AOI22M1P U216 ( .A(n45), .B(\Queue[2][14] ), .C(\Queue[1][14] ), .D(n42), 
        .Z(n80) );
  OAI21M1P U217 ( .A(n47), .B(n180), .C(n80), .Z(n435) );
  AOI22M1P U218 ( .A(n46), .B(\Queue[2][15] ), .C(\Queue[1][15] ), .D(n42), 
        .Z(n81) );
  OAI21M1P U219 ( .A(n47), .B(n182), .C(n81), .Z(n436) );
  AOI22M1P U220 ( .A(n45), .B(\Queue[2][16] ), .C(\Queue[1][16] ), .D(n42), 
        .Z(n82) );
  OAI21M1P U221 ( .A(n47), .B(n184), .C(n82), .Z(n437) );
  AOI22M1P U222 ( .A(n46), .B(\Queue[2][17] ), .C(\Queue[1][17] ), .D(n42), 
        .Z(n83) );
  OAI21M1P U223 ( .A(n47), .B(n186), .C(n83), .Z(n438) );
  AOI22M1P U224 ( .A(n45), .B(\Queue[2][18] ), .C(\Queue[1][18] ), .D(n43), 
        .Z(n84) );
  OAI21M1P U225 ( .A(n47), .B(n188), .C(n84), .Z(n439) );
  AOI22M1P U226 ( .A(n46), .B(\Queue[2][19] ), .C(\Queue[1][19] ), .D(n43), 
        .Z(n85) );
  OAI21M1P U227 ( .A(n47), .B(n190), .C(n85), .Z(n440) );
  AOI22M1P U228 ( .A(n46), .B(\Queue[2][20] ), .C(\Queue[1][20] ), .D(n43), 
        .Z(n86) );
  OAI21M1P U229 ( .A(n47), .B(n192), .C(n86), .Z(n441) );
  AOI22M1P U230 ( .A(n45), .B(\Queue[2][21] ), .C(\Queue[1][21] ), .D(n43), 
        .Z(n87) );
  OAI21M1P U231 ( .A(n47), .B(n194), .C(n87), .Z(n442) );
  AOI22M1P U232 ( .A(n45), .B(\Queue[2][22] ), .C(\Queue[1][22] ), .D(n43), 
        .Z(n88) );
  OAI21M1P U233 ( .A(n47), .B(n196), .C(n88), .Z(n443) );
  AOI22M1P U234 ( .A(n45), .B(\Queue[2][23] ), .C(\Queue[1][23] ), .D(n43), 
        .Z(n89) );
  OAI21M1P U235 ( .A(n47), .B(n198), .C(n89), .Z(n444) );
  AOI22M1P U236 ( .A(n45), .B(\Queue[2][24] ), .C(\Queue[1][24] ), .D(n43), 
        .Z(n90) );
  OAI21M1P U237 ( .A(n47), .B(n200), .C(n90), .Z(n445) );
  AOI22M1P U238 ( .A(n45), .B(\Queue[2][25] ), .C(\Queue[1][25] ), .D(n43), 
        .Z(n91) );
  OAI21M1P U239 ( .A(n47), .B(n202), .C(n91), .Z(n446) );
  AOI22M1P U240 ( .A(n45), .B(\Queue[2][26] ), .C(\Queue[1][26] ), .D(n43), 
        .Z(n92) );
  OAI21M1P U241 ( .A(n47), .B(n204), .C(n92), .Z(n447) );
  AOI22M1P U242 ( .A(n45), .B(\Queue[2][27] ), .C(\Queue[1][27] ), .D(n44), 
        .Z(n93) );
  OAI21M1P U243 ( .A(n47), .B(n206), .C(n93), .Z(n448) );
  AOI22M1P U244 ( .A(n45), .B(\Queue[2][28] ), .C(\Queue[1][28] ), .D(n44), 
        .Z(n94) );
  OAI21M1P U245 ( .A(n47), .B(n208), .C(n94), .Z(n449) );
  AOI22M1P U246 ( .A(n45), .B(\Queue[2][29] ), .C(\Queue[1][29] ), .D(n44), 
        .Z(n95) );
  OAI21M1P U247 ( .A(n47), .B(n374), .C(n95), .Z(n450) );
  AOI22M1P U248 ( .A(n45), .B(\Queue[2][30] ), .C(\Queue[1][30] ), .D(n44), 
        .Z(n96) );
  OAI21M1P U249 ( .A(n47), .B(n376), .C(n96), .Z(n451) );
  AOI22M1P U250 ( .A(n45), .B(\Queue[2][31] ), .C(\Queue[1][31] ), .D(n44), 
        .Z(n99) );
  OAI21M1P U251 ( .A(n47), .B(n381), .C(n99), .Z(n452) );
  AOI22M1P U252 ( .A(\Queue[1][0] ), .B(n136), .C(n135), .D(Packet_Out[0]), 
        .Z(n104) );
  OAI21M1P U253 ( .A(n152), .B(n4), .C(n104), .Z(n453) );
  AOI22M1P U254 ( .A(\Queue[1][1] ), .B(n136), .C(n135), .D(Packet_Out[1]), 
        .Z(n105) );
  OAI21M1P U255 ( .A(n154), .B(n4), .C(n105), .Z(n454) );
  AOI22M1P U256 ( .A(\Queue[1][2] ), .B(n136), .C(n135), .D(Packet_Out[2]), 
        .Z(n106) );
  OAI21M1P U257 ( .A(n156), .B(n4), .C(n106), .Z(n455) );
  AOI22M1P U258 ( .A(\Queue[1][3] ), .B(n136), .C(n135), .D(Packet_Out[3]), 
        .Z(n107) );
  OAI21M1P U259 ( .A(n158), .B(n4), .C(n107), .Z(n456) );
  AOI22M1P U260 ( .A(\Queue[1][4] ), .B(n136), .C(n135), .D(Packet_Out[4]), 
        .Z(n108) );
  OAI21M1P U261 ( .A(n160), .B(n4), .C(n108), .Z(n457) );
  AOI22M1P U262 ( .A(\Queue[1][5] ), .B(n136), .C(n135), .D(Packet_Out[5]), 
        .Z(n109) );
  OAI21M1P U263 ( .A(n162), .B(n4), .C(n109), .Z(n458) );
  AOI22M1P U264 ( .A(\Queue[1][6] ), .B(n136), .C(n135), .D(Packet_Out[6]), 
        .Z(n110) );
  OAI21M1P U265 ( .A(n164), .B(n4), .C(n110), .Z(n459) );
  AOI22M1P U266 ( .A(\Queue[1][7] ), .B(n136), .C(n135), .D(Packet_Out[7]), 
        .Z(n111) );
  OAI21M1P U267 ( .A(n166), .B(n4), .C(n111), .Z(n460) );
  AOI22M1P U268 ( .A(\Queue[1][8] ), .B(n136), .C(n135), .D(Packet_Out[8]), 
        .Z(n112) );
  OAI21M1P U269 ( .A(n168), .B(n4), .C(n112), .Z(n461) );
  AOI22M1P U270 ( .A(\Queue[1][9] ), .B(n136), .C(n135), .D(Packet_Out[9]), 
        .Z(n113) );
  OAI21M1P U271 ( .A(n170), .B(n4), .C(n113), .Z(n462) );
  AOI22M1P U272 ( .A(\Queue[1][10] ), .B(n136), .C(n135), .D(Packet_Out[10]), 
        .Z(n114) );
  OAI21M1P U273 ( .A(n172), .B(n4), .C(n114), .Z(n463) );
  AOI22M1P U274 ( .A(\Queue[1][11] ), .B(n136), .C(n135), .D(Packet_Out[11]), 
        .Z(n115) );
  OAI21M1P U275 ( .A(n174), .B(n4), .C(n115), .Z(n464) );
  AOI22M1P U276 ( .A(\Queue[1][12] ), .B(n136), .C(n135), .D(Packet_Out[12]), 
        .Z(n116) );
  OAI21M1P U277 ( .A(n176), .B(n4), .C(n116), .Z(n465) );
  AOI22M1P U278 ( .A(\Queue[1][13] ), .B(n136), .C(n135), .D(Packet_Out[13]), 
        .Z(n117) );
  OAI21M1P U279 ( .A(n178), .B(n4), .C(n117), .Z(n466) );
  AOI22M1P U280 ( .A(\Queue[1][14] ), .B(n136), .C(n135), .D(Packet_Out[14]), 
        .Z(n118) );
  OAI21M1P U281 ( .A(n180), .B(n4), .C(n118), .Z(n467) );
  AOI22M1P U282 ( .A(\Queue[1][15] ), .B(n136), .C(n135), .D(Packet_Out[15]), 
        .Z(n119) );
  OAI21M1P U283 ( .A(n182), .B(n4), .C(n119), .Z(n468) );
  AOI22M1P U284 ( .A(\Queue[1][16] ), .B(n136), .C(n135), .D(Packet_Out[16]), 
        .Z(n120) );
  OAI21M1P U285 ( .A(n184), .B(n4), .C(n120), .Z(n469) );
  AOI22M1P U286 ( .A(\Queue[1][17] ), .B(n136), .C(n135), .D(Packet_Out[17]), 
        .Z(n121) );
  OAI21M1P U287 ( .A(n186), .B(n4), .C(n121), .Z(n470) );
  AOI22M1P U288 ( .A(\Queue[1][18] ), .B(n136), .C(n135), .D(Packet_Out[18]), 
        .Z(n122) );
  OAI21M1P U289 ( .A(n188), .B(n4), .C(n122), .Z(n471) );
  AOI22M1P U290 ( .A(\Queue[1][19] ), .B(n136), .C(n135), .D(Packet_Out[19]), 
        .Z(n123) );
  OAI21M1P U291 ( .A(n190), .B(n4), .C(n123), .Z(n472) );
  AOI22M1P U292 ( .A(\Queue[1][20] ), .B(n136), .C(n135), .D(Packet_Out[20]), 
        .Z(n124) );
  OAI21M1P U293 ( .A(n192), .B(n4), .C(n124), .Z(n473) );
  AOI22M1P U294 ( .A(\Queue[1][21] ), .B(n136), .C(n135), .D(Packet_Out[21]), 
        .Z(n125) );
  OAI21M1P U295 ( .A(n194), .B(n4), .C(n125), .Z(n474) );
  AOI22M1P U296 ( .A(\Queue[1][22] ), .B(n136), .C(n135), .D(Packet_Out[22]), 
        .Z(n126) );
  OAI21M1P U297 ( .A(n196), .B(n4), .C(n126), .Z(n475) );
  AOI22M1P U298 ( .A(\Queue[1][23] ), .B(n136), .C(n135), .D(Packet_Out[23]), 
        .Z(n127) );
  OAI21M1P U299 ( .A(n198), .B(n4), .C(n127), .Z(n476) );
  AOI22M1P U300 ( .A(\Queue[1][24] ), .B(n136), .C(n135), .D(Packet_Out[24]), 
        .Z(n128) );
  OAI21M1P U301 ( .A(n200), .B(n4), .C(n128), .Z(n477) );
  AOI22M1P U302 ( .A(\Queue[1][25] ), .B(n136), .C(n135), .D(Packet_Out[25]), 
        .Z(n129) );
  OAI21M1P U303 ( .A(n202), .B(n4), .C(n129), .Z(n478) );
  AOI22M1P U304 ( .A(\Queue[1][26] ), .B(n136), .C(n135), .D(Packet_Out[26]), 
        .Z(n130) );
  OAI21M1P U305 ( .A(n204), .B(n4), .C(n130), .Z(n479) );
  AOI22M1P U306 ( .A(\Queue[1][27] ), .B(n136), .C(n135), .D(Packet_Out[27]), 
        .Z(n131) );
  OAI21M1P U307 ( .A(n206), .B(n4), .C(n131), .Z(n480) );
  AOI22M1P U308 ( .A(\Queue[1][28] ), .B(n136), .C(n135), .D(Packet_Out[28]), 
        .Z(n132) );
  OAI21M1P U309 ( .A(n208), .B(n4), .C(n132), .Z(n481) );
  AOI22M1P U310 ( .A(\Queue[1][29] ), .B(n136), .C(n135), .D(Packet_Out[29]), 
        .Z(n133) );
  OAI21M1P U311 ( .A(n374), .B(n4), .C(n133), .Z(n482) );
  AOI22M1P U312 ( .A(\Queue[1][30] ), .B(n136), .C(n135), .D(Packet_Out[30]), 
        .Z(n134) );
  OAI21M1P U313 ( .A(n376), .B(n4), .C(n134), .Z(n483) );
  AOI22M1P U314 ( .A(\Queue[1][31] ), .B(n136), .C(n135), .D(Packet_Out[31]), 
        .Z(n137) );
  OAI21M1P U315 ( .A(n381), .B(n4), .C(n137), .Z(n484) );
  ND2M1P U316 ( .A(n139), .B(n146), .Z(n147) );
  AOI21M1P U317 ( .A(Write_Ack), .B(n149), .C(n150), .Z(n143) );
  AOI22M1P U318 ( .A(\Queue[2][0] ), .B(n51), .C(\Queue[3][0] ), .D(n50), .Z(
        n141) );
  AOI22M1P U319 ( .A(\Queue[2][30] ), .B(n51), .C(n49), .D(\Queue[3][30] ), 
        .Z(n142) );
  OAI21M1P U320 ( .A(n376), .B(n52), .C(n142), .Z(n515) );
  AOI22M1P U321 ( .A(\Queue[2][31] ), .B(n51), .C(n49), .D(\Queue[3][31] ), 
        .Z(n145) );
  OAI21M1P U322 ( .A(n381), .B(n52), .C(n145), .Z(n516) );
  AOI22M1P U323 ( .A(\Queue[3][1] ), .B(n53), .C(n377), .D(\Queue[4][1] ), .Z(
        n153) );
  OAI21M1P U324 ( .A(n154), .B(n380), .C(n153), .Z(n518) );
  AOI22M1P U325 ( .A(\Queue[3][2] ), .B(n53), .C(n377), .D(\Queue[4][2] ), .Z(
        n155) );
  OAI21M1P U326 ( .A(n156), .B(n380), .C(n155), .Z(n519) );
  AOI22M1P U327 ( .A(\Queue[3][3] ), .B(n53), .C(n377), .D(\Queue[4][3] ), .Z(
        n157) );
  OAI21M1P U328 ( .A(n158), .B(n380), .C(n157), .Z(n520) );
  AOI22M1P U329 ( .A(\Queue[3][4] ), .B(n53), .C(n377), .D(\Queue[4][4] ), .Z(
        n159) );
  OAI21M1P U330 ( .A(n160), .B(n380), .C(n159), .Z(n521) );
  AOI22M1P U331 ( .A(\Queue[3][5] ), .B(n53), .C(n377), .D(\Queue[4][5] ), .Z(
        n161) );
  OAI21M1P U332 ( .A(n162), .B(n380), .C(n161), .Z(n522) );
  AOI22M1P U333 ( .A(\Queue[3][6] ), .B(n53), .C(n377), .D(\Queue[4][6] ), .Z(
        n163) );
  OAI21M1P U334 ( .A(n164), .B(n380), .C(n163), .Z(n523) );
  AOI22M1P U335 ( .A(\Queue[3][7] ), .B(n53), .C(n377), .D(\Queue[4][7] ), .Z(
        n165) );
  OAI21M1P U336 ( .A(n166), .B(n380), .C(n165), .Z(n524) );
  AOI22M1P U337 ( .A(\Queue[3][8] ), .B(n53), .C(n377), .D(\Queue[4][8] ), .Z(
        n167) );
  OAI21M1P U338 ( .A(n168), .B(n380), .C(n167), .Z(n525) );
  AOI22M1P U339 ( .A(\Queue[3][9] ), .B(n53), .C(n377), .D(\Queue[4][9] ), .Z(
        n169) );
  OAI21M1P U340 ( .A(n170), .B(n380), .C(n169), .Z(n526) );
  AOI22M1P U341 ( .A(\Queue[3][10] ), .B(n53), .C(n377), .D(\Queue[4][10] ), 
        .Z(n171) );
  OAI21M1P U342 ( .A(n172), .B(n380), .C(n171), .Z(n527) );
  AOI22M1P U343 ( .A(\Queue[3][11] ), .B(n53), .C(n377), .D(\Queue[4][11] ), 
        .Z(n173) );
  OAI21M1P U344 ( .A(n174), .B(n380), .C(n173), .Z(n528) );
  AOI22M1P U345 ( .A(\Queue[3][12] ), .B(n53), .C(n377), .D(\Queue[4][12] ), 
        .Z(n175) );
  OAI21M1P U346 ( .A(n176), .B(n380), .C(n175), .Z(n529) );
  AOI22M1P U347 ( .A(\Queue[3][13] ), .B(n53), .C(n377), .D(\Queue[4][13] ), 
        .Z(n177) );
  OAI21M1P U348 ( .A(n178), .B(n380), .C(n177), .Z(n530) );
  AOI22M1P U349 ( .A(\Queue[3][14] ), .B(n53), .C(n377), .D(\Queue[4][14] ), 
        .Z(n179) );
  OAI21M1P U350 ( .A(n180), .B(n380), .C(n179), .Z(n531) );
  AOI22M1P U351 ( .A(\Queue[3][15] ), .B(n53), .C(n377), .D(\Queue[4][15] ), 
        .Z(n181) );
  OAI21M1P U352 ( .A(n182), .B(n380), .C(n181), .Z(n532) );
  AOI22M1P U353 ( .A(\Queue[3][16] ), .B(n53), .C(n377), .D(\Queue[4][16] ), 
        .Z(n183) );
  OAI21M1P U354 ( .A(n184), .B(n380), .C(n183), .Z(n533) );
  AOI22M1P U355 ( .A(\Queue[3][17] ), .B(n53), .C(n377), .D(\Queue[4][17] ), 
        .Z(n185) );
  OAI21M1P U356 ( .A(n186), .B(n380), .C(n185), .Z(n534) );
  AOI22M1P U357 ( .A(\Queue[3][18] ), .B(n53), .C(n377), .D(\Queue[4][18] ), 
        .Z(n187) );
  OAI21M1P U358 ( .A(n188), .B(n380), .C(n187), .Z(n535) );
  AOI22M1P U359 ( .A(\Queue[3][19] ), .B(n53), .C(n377), .D(\Queue[4][19] ), 
        .Z(n189) );
  OAI21M1P U360 ( .A(n190), .B(n380), .C(n189), .Z(n536) );
  AOI22M1P U361 ( .A(\Queue[3][20] ), .B(n378), .C(n377), .D(\Queue[4][20] ), 
        .Z(n191) );
  OAI21M1P U362 ( .A(n192), .B(n380), .C(n191), .Z(n537) );
  AOI22M1P U363 ( .A(\Queue[3][21] ), .B(n378), .C(n377), .D(\Queue[4][21] ), 
        .Z(n193) );
  OAI21M1P U364 ( .A(n194), .B(n380), .C(n193), .Z(n538) );
  AOI22M1P U365 ( .A(\Queue[3][22] ), .B(n378), .C(n377), .D(\Queue[4][22] ), 
        .Z(n195) );
  OAI21M1P U366 ( .A(n196), .B(n380), .C(n195), .Z(n539) );
  AOI22M1P U367 ( .A(\Queue[3][23] ), .B(n53), .C(n377), .D(\Queue[4][23] ), 
        .Z(n197) );
  OAI21M1P U368 ( .A(n198), .B(n380), .C(n197), .Z(n540) );
  AOI22M1P U369 ( .A(\Queue[3][24] ), .B(n53), .C(n377), .D(\Queue[4][24] ), 
        .Z(n199) );
  OAI21M1P U370 ( .A(n200), .B(n380), .C(n199), .Z(n541) );
  AOI22M1P U371 ( .A(\Queue[3][25] ), .B(n53), .C(n377), .D(\Queue[4][25] ), 
        .Z(n201) );
  OAI21M1P U372 ( .A(n202), .B(n380), .C(n201), .Z(n542) );
  AOI22M1P U373 ( .A(\Queue[3][26] ), .B(n53), .C(n377), .D(\Queue[4][26] ), 
        .Z(n203) );
  OAI21M1P U374 ( .A(n204), .B(n380), .C(n203), .Z(n543) );
  AOI22M1P U375 ( .A(\Queue[3][27] ), .B(n53), .C(n377), .D(\Queue[4][27] ), 
        .Z(n205) );
  OAI21M1P U376 ( .A(n206), .B(n380), .C(n205), .Z(n544) );
  AOI22M1P U377 ( .A(\Queue[3][28] ), .B(n53), .C(n377), .D(\Queue[4][28] ), 
        .Z(n207) );
  OAI21M1P U378 ( .A(n208), .B(n380), .C(n207), .Z(n545) );
  AOI22M1P U379 ( .A(\Queue[3][29] ), .B(n53), .C(n377), .D(\Queue[4][29] ), 
        .Z(n373) );
  OAI21M1P U380 ( .A(n374), .B(n380), .C(n373), .Z(n546) );
  AOI22M1P U381 ( .A(\Queue[3][30] ), .B(n53), .C(n377), .D(\Queue[4][30] ), 
        .Z(n375) );
  OAI21M1P U382 ( .A(n376), .B(n380), .C(n375), .Z(n547) );
  AOI22M1P U383 ( .A(\Queue[3][31] ), .B(n53), .C(n377), .D(\Queue[4][31] ), 
        .Z(n379) );
  OAI21M1P U384 ( .A(n381), .B(n380), .C(n379), .Z(n548) );
  N1M1P U385 ( .A(n549), .Z(Empty) );
  AOI22M1P U386 ( .A(n384), .B(n383), .C(n382), .D(Empty), .Z(n550) );
endmodule


module Packet_Queue_8 ( Clk_r, Rst_n, Packet_In, Read_Ack, Write_Ack, 
        Packet_Out, Empty, Full );
  input [31:0] Packet_In;
  output [31:0] Packet_Out;
  input Clk_r, Rst_n, Read_Ack, Write_Ack;
  output Empty, Full;
  wire   \Queue[4][31] , \Queue[4][30] , \Queue[4][29] , \Queue[4][28] ,
         \Queue[4][27] , \Queue[4][26] , \Queue[4][25] , \Queue[4][24] ,
         \Queue[4][23] , \Queue[4][22] , \Queue[4][21] , \Queue[4][20] ,
         \Queue[4][19] , \Queue[4][18] , \Queue[4][17] , \Queue[4][16] ,
         \Queue[4][15] , \Queue[4][14] , \Queue[4][13] , \Queue[4][12] ,
         \Queue[4][11] , \Queue[4][10] , \Queue[4][9] , \Queue[4][8] ,
         \Queue[4][7] , \Queue[4][6] , \Queue[4][5] , \Queue[4][4] ,
         \Queue[4][3] , \Queue[4][2] , \Queue[4][1] , \Queue[4][0] ,
         \Queue[3][31] , \Queue[3][30] , \Queue[3][29] , \Queue[3][28] ,
         \Queue[3][27] , \Queue[3][26] , \Queue[3][25] , \Queue[3][24] ,
         \Queue[3][23] , \Queue[3][22] , \Queue[3][21] , \Queue[3][20] ,
         \Queue[3][19] , \Queue[3][18] , \Queue[3][17] , \Queue[3][16] ,
         \Queue[3][15] , \Queue[3][14] , \Queue[3][13] , \Queue[3][12] ,
         \Queue[3][11] , \Queue[3][10] , \Queue[3][9] , \Queue[3][8] ,
         \Queue[3][7] , \Queue[3][6] , \Queue[3][5] , \Queue[3][4] ,
         \Queue[3][3] , \Queue[3][2] , \Queue[3][1] , \Queue[3][0] ,
         \Queue[2][31] , \Queue[2][30] , \Queue[2][29] , \Queue[2][28] ,
         \Queue[2][27] , \Queue[2][26] , \Queue[2][25] , \Queue[2][24] ,
         \Queue[2][23] , \Queue[2][22] , \Queue[2][21] , \Queue[2][20] ,
         \Queue[2][19] , \Queue[2][18] , \Queue[2][17] , \Queue[2][16] ,
         \Queue[2][15] , \Queue[2][14] , \Queue[2][13] , \Queue[2][12] ,
         \Queue[2][11] , \Queue[2][10] , \Queue[2][9] , \Queue[2][8] ,
         \Queue[2][7] , \Queue[2][6] , \Queue[2][5] , \Queue[2][4] ,
         \Queue[2][3] , \Queue[2][2] , \Queue[2][1] , \Queue[2][0] ,
         \Queue[1][31] , \Queue[1][30] , \Queue[1][29] , \Queue[1][28] ,
         \Queue[1][27] , \Queue[1][26] , \Queue[1][25] , \Queue[1][24] ,
         \Queue[1][23] , \Queue[1][22] , \Queue[1][21] , \Queue[1][20] ,
         \Queue[1][19] , \Queue[1][18] , \Queue[1][17] , \Queue[1][16] ,
         \Queue[1][15] , \Queue[1][14] , \Queue[1][13] , \Queue[1][12] ,
         \Queue[1][11] , \Queue[1][10] , \Queue[1][9] , \Queue[1][8] ,
         \Queue[1][7] , \Queue[1][6] , \Queue[1][5] , \Queue[1][4] ,
         \Queue[1][3] , \Queue[1][2] , \Queue[1][1] , \Queue[1][0] , n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542;
  wire   [2:0] Count;

  FDN2QM1P \Count_reg[0]  ( .D(n377), .CPN(Clk_r), .CD(Rst_n), .Q(Count[0]) );
  FDN2QM1P \Count_reg[1]  ( .D(n378), .CPN(Clk_r), .CD(Rst_n), .Q(Count[1]) );
  FDN2QM1P \Count_reg[2]  ( .D(n379), .CPN(Clk_r), .CD(Rst_n), .Q(Count[2]) );
  FDN1QM1P \Queue_reg[4][30]  ( .D(n411), .CPN(Clk_r), .Q(\Queue[4][30] ) );
  FDN1QM1P \Queue_reg[3][30]  ( .D(n539), .CPN(Clk_r), .Q(\Queue[3][30] ) );
  FDN1QM1P \Queue_reg[2][30]  ( .D(n507), .CPN(Clk_r), .Q(\Queue[2][30] ) );
  FDN1QM1P \Queue_reg[4][29]  ( .D(n410), .CPN(Clk_r), .Q(\Queue[4][29] ) );
  FDN1QM1P \Queue_reg[3][29]  ( .D(n538), .CPN(Clk_r), .Q(\Queue[3][29] ) );
  FDN1QM1P \Queue_reg[2][29]  ( .D(n506), .CPN(Clk_r), .Q(\Queue[2][29] ) );
  FDN1QM1P \Queue_reg[4][28]  ( .D(n409), .CPN(Clk_r), .Q(\Queue[4][28] ) );
  FDN1QM1P \Queue_reg[3][28]  ( .D(n537), .CPN(Clk_r), .Q(\Queue[3][28] ) );
  FDN1QM1P \Queue_reg[2][28]  ( .D(n505), .CPN(Clk_r), .Q(\Queue[2][28] ) );
  FDN1QM1P \Queue_reg[4][27]  ( .D(n408), .CPN(Clk_r), .Q(\Queue[4][27] ) );
  FDN1QM1P \Queue_reg[3][27]  ( .D(n536), .CPN(Clk_r), .Q(\Queue[3][27] ) );
  FDN1QM1P \Queue_reg[2][27]  ( .D(n504), .CPN(Clk_r), .Q(\Queue[2][27] ) );
  FDN1QM1P \Queue_reg[4][26]  ( .D(n407), .CPN(Clk_r), .Q(\Queue[4][26] ) );
  FDN1QM1P \Queue_reg[3][26]  ( .D(n535), .CPN(Clk_r), .Q(\Queue[3][26] ) );
  FDN1QM1P \Queue_reg[2][26]  ( .D(n503), .CPN(Clk_r), .Q(\Queue[2][26] ) );
  FDN1QM1P \Queue_reg[4][25]  ( .D(n406), .CPN(Clk_r), .Q(\Queue[4][25] ) );
  FDN1QM1P \Queue_reg[3][25]  ( .D(n534), .CPN(Clk_r), .Q(\Queue[3][25] ) );
  FDN1QM1P \Queue_reg[2][25]  ( .D(n502), .CPN(Clk_r), .Q(\Queue[2][25] ) );
  FDN1QM1P \Queue_reg[4][24]  ( .D(n405), .CPN(Clk_r), .Q(\Queue[4][24] ) );
  FDN1QM1P \Queue_reg[3][24]  ( .D(n533), .CPN(Clk_r), .Q(\Queue[3][24] ) );
  FDN1QM1P \Queue_reg[2][24]  ( .D(n501), .CPN(Clk_r), .Q(\Queue[2][24] ) );
  FDN1QM1P \Queue_reg[4][23]  ( .D(n404), .CPN(Clk_r), .Q(\Queue[4][23] ) );
  FDN1QM1P \Queue_reg[3][23]  ( .D(n532), .CPN(Clk_r), .Q(\Queue[3][23] ) );
  FDN1QM1P \Queue_reg[2][23]  ( .D(n500), .CPN(Clk_r), .Q(\Queue[2][23] ) );
  FDN1QM1P \Queue_reg[4][22]  ( .D(n403), .CPN(Clk_r), .Q(\Queue[4][22] ) );
  FDN1QM1P \Queue_reg[3][22]  ( .D(n531), .CPN(Clk_r), .Q(\Queue[3][22] ) );
  FDN1QM1P \Queue_reg[2][22]  ( .D(n499), .CPN(Clk_r), .Q(\Queue[2][22] ) );
  FDN1QM1P \Queue_reg[4][21]  ( .D(n402), .CPN(Clk_r), .Q(\Queue[4][21] ) );
  FDN1QM1P \Queue_reg[3][21]  ( .D(n530), .CPN(Clk_r), .Q(\Queue[3][21] ) );
  FDN1QM1P \Queue_reg[2][21]  ( .D(n498), .CPN(Clk_r), .Q(\Queue[2][21] ) );
  FDN1QM1P \Queue_reg[4][20]  ( .D(n401), .CPN(Clk_r), .Q(\Queue[4][20] ) );
  FDN1QM1P \Queue_reg[3][20]  ( .D(n529), .CPN(Clk_r), .Q(\Queue[3][20] ) );
  FDN1QM1P \Queue_reg[2][20]  ( .D(n497), .CPN(Clk_r), .Q(\Queue[2][20] ) );
  FDN1QM1P \Queue_reg[4][19]  ( .D(n400), .CPN(Clk_r), .Q(\Queue[4][19] ) );
  FDN1QM1P \Queue_reg[3][19]  ( .D(n528), .CPN(Clk_r), .Q(\Queue[3][19] ) );
  FDN1QM1P \Queue_reg[2][19]  ( .D(n496), .CPN(Clk_r), .Q(\Queue[2][19] ) );
  FDN1QM1P \Queue_reg[4][18]  ( .D(n399), .CPN(Clk_r), .Q(\Queue[4][18] ) );
  FDN1QM1P \Queue_reg[3][18]  ( .D(n527), .CPN(Clk_r), .Q(\Queue[3][18] ) );
  FDN1QM1P \Queue_reg[2][18]  ( .D(n495), .CPN(Clk_r), .Q(\Queue[2][18] ) );
  FDN1QM1P \Queue_reg[4][17]  ( .D(n398), .CPN(Clk_r), .Q(\Queue[4][17] ) );
  FDN1QM1P \Queue_reg[3][17]  ( .D(n526), .CPN(Clk_r), .Q(\Queue[3][17] ) );
  FDN1QM1P \Queue_reg[2][17]  ( .D(n494), .CPN(Clk_r), .Q(\Queue[2][17] ) );
  FDN1QM1P \Queue_reg[4][16]  ( .D(n397), .CPN(Clk_r), .Q(\Queue[4][16] ) );
  FDN1QM1P \Queue_reg[3][16]  ( .D(n525), .CPN(Clk_r), .Q(\Queue[3][16] ) );
  FDN1QM1P \Queue_reg[2][16]  ( .D(n493), .CPN(Clk_r), .Q(\Queue[2][16] ) );
  FDN1QM1P \Queue_reg[4][15]  ( .D(n396), .CPN(Clk_r), .Q(\Queue[4][15] ) );
  FDN1QM1P \Queue_reg[3][15]  ( .D(n524), .CPN(Clk_r), .Q(\Queue[3][15] ) );
  FDN1QM1P \Queue_reg[2][15]  ( .D(n492), .CPN(Clk_r), .Q(\Queue[2][15] ) );
  FDN1QM1P \Queue_reg[4][14]  ( .D(n395), .CPN(Clk_r), .Q(\Queue[4][14] ) );
  FDN1QM1P \Queue_reg[3][14]  ( .D(n523), .CPN(Clk_r), .Q(\Queue[3][14] ) );
  FDN1QM1P \Queue_reg[2][14]  ( .D(n491), .CPN(Clk_r), .Q(\Queue[2][14] ) );
  FDN1QM1P \Queue_reg[4][13]  ( .D(n394), .CPN(Clk_r), .Q(\Queue[4][13] ) );
  FDN1QM1P \Queue_reg[3][13]  ( .D(n522), .CPN(Clk_r), .Q(\Queue[3][13] ) );
  FDN1QM1P \Queue_reg[2][13]  ( .D(n490), .CPN(Clk_r), .Q(\Queue[2][13] ) );
  FDN1QM1P \Queue_reg[4][12]  ( .D(n393), .CPN(Clk_r), .Q(\Queue[4][12] ) );
  FDN1QM1P \Queue_reg[3][12]  ( .D(n521), .CPN(Clk_r), .Q(\Queue[3][12] ) );
  FDN1QM1P \Queue_reg[2][12]  ( .D(n489), .CPN(Clk_r), .Q(\Queue[2][12] ) );
  FDN1QM1P \Queue_reg[4][11]  ( .D(n392), .CPN(Clk_r), .Q(\Queue[4][11] ) );
  FDN1QM1P \Queue_reg[3][11]  ( .D(n520), .CPN(Clk_r), .Q(\Queue[3][11] ) );
  FDN1QM1P \Queue_reg[2][11]  ( .D(n488), .CPN(Clk_r), .Q(\Queue[2][11] ) );
  FDN1QM1P \Queue_reg[4][10]  ( .D(n391), .CPN(Clk_r), .Q(\Queue[4][10] ) );
  FDN1QM1P \Queue_reg[3][10]  ( .D(n519), .CPN(Clk_r), .Q(\Queue[3][10] ) );
  FDN1QM1P \Queue_reg[2][10]  ( .D(n487), .CPN(Clk_r), .Q(\Queue[2][10] ) );
  FDN1QM1P \Queue_reg[4][9]  ( .D(n390), .CPN(Clk_r), .Q(\Queue[4][9] ) );
  FDN1QM1P \Queue_reg[3][9]  ( .D(n518), .CPN(Clk_r), .Q(\Queue[3][9] ) );
  FDN1QM1P \Queue_reg[2][9]  ( .D(n486), .CPN(Clk_r), .Q(\Queue[2][9] ) );
  FDN1QM1P \Queue_reg[4][8]  ( .D(n389), .CPN(Clk_r), .Q(\Queue[4][8] ) );
  FDN1QM1P \Queue_reg[3][8]  ( .D(n517), .CPN(Clk_r), .Q(\Queue[3][8] ) );
  FDN1QM1P \Queue_reg[2][8]  ( .D(n485), .CPN(Clk_r), .Q(\Queue[2][8] ) );
  FDN1QM1P \Queue_reg[4][7]  ( .D(n388), .CPN(Clk_r), .Q(\Queue[4][7] ) );
  FDN1QM1P \Queue_reg[3][7]  ( .D(n516), .CPN(Clk_r), .Q(\Queue[3][7] ) );
  FDN1QM1P \Queue_reg[2][7]  ( .D(n484), .CPN(Clk_r), .Q(\Queue[2][7] ) );
  FDN1QM1P \Queue_reg[4][6]  ( .D(n387), .CPN(Clk_r), .Q(\Queue[4][6] ) );
  FDN1QM1P \Queue_reg[3][6]  ( .D(n515), .CPN(Clk_r), .Q(\Queue[3][6] ) );
  FDN1QM1P \Queue_reg[2][6]  ( .D(n483), .CPN(Clk_r), .Q(\Queue[2][6] ) );
  FDN1QM1P \Queue_reg[4][5]  ( .D(n386), .CPN(Clk_r), .Q(\Queue[4][5] ) );
  FDN1QM1P \Queue_reg[3][5]  ( .D(n514), .CPN(Clk_r), .Q(\Queue[3][5] ) );
  FDN1QM1P \Queue_reg[2][5]  ( .D(n482), .CPN(Clk_r), .Q(\Queue[2][5] ) );
  FDN1QM1P \Queue_reg[4][4]  ( .D(n385), .CPN(Clk_r), .Q(\Queue[4][4] ) );
  FDN1QM1P \Queue_reg[3][4]  ( .D(n513), .CPN(Clk_r), .Q(\Queue[3][4] ) );
  FDN1QM1P \Queue_reg[2][4]  ( .D(n481), .CPN(Clk_r), .Q(\Queue[2][4] ) );
  FDN1QM1P \Queue_reg[4][3]  ( .D(n384), .CPN(Clk_r), .Q(\Queue[4][3] ) );
  FDN1QM1P \Queue_reg[3][3]  ( .D(n512), .CPN(Clk_r), .Q(\Queue[3][3] ) );
  FDN1QM1P \Queue_reg[2][3]  ( .D(n480), .CPN(Clk_r), .Q(\Queue[2][3] ) );
  FDN1QM1P \Queue_reg[4][2]  ( .D(n383), .CPN(Clk_r), .Q(\Queue[4][2] ) );
  FDN1QM1P \Queue_reg[3][2]  ( .D(n511), .CPN(Clk_r), .Q(\Queue[3][2] ) );
  FDN1QM1P \Queue_reg[2][2]  ( .D(n479), .CPN(Clk_r), .Q(\Queue[2][2] ) );
  FDN1QM1P \Queue_reg[4][1]  ( .D(n382), .CPN(Clk_r), .Q(\Queue[4][1] ) );
  FDN1QM1P \Queue_reg[3][1]  ( .D(n510), .CPN(Clk_r), .Q(\Queue[3][1] ) );
  FDN1QM1P \Queue_reg[2][1]  ( .D(n478), .CPN(Clk_r), .Q(\Queue[2][1] ) );
  FDN1QM1P \Queue_reg[4][0]  ( .D(n381), .CPN(Clk_r), .Q(\Queue[4][0] ) );
  FDN1QM1P \Queue_reg[3][0]  ( .D(n509), .CPN(Clk_r), .Q(\Queue[3][0] ) );
  FDN1QM1P \Queue_reg[2][0]  ( .D(n477), .CPN(Clk_r), .Q(\Queue[2][0] ) );
  FDN1QM1P \Queue_reg[4][31]  ( .D(n380), .CPN(Clk_r), .Q(\Queue[4][31] ) );
  FDN1QM1P \Queue_reg[3][31]  ( .D(n540), .CPN(Clk_r), .Q(\Queue[3][31] ) );
  FDN1QM1P \Queue_reg[2][31]  ( .D(n508), .CPN(Clk_r), .Q(\Queue[2][31] ) );
  FDN2QM1P Full_reg ( .D(n412), .CPN(Clk_r), .CD(Rst_n), .Q(Full) );
  FDN1QM1P \Queue_reg[1][31]  ( .D(n444), .CPN(Clk_r), .Q(\Queue[1][31] ) );
  FDN1QM1P \Queue_reg[0][31]  ( .D(n476), .CPN(Clk_r), .Q(Packet_Out[31]) );
  FDN1QM1P \Queue_reg[1][30]  ( .D(n443), .CPN(Clk_r), .Q(\Queue[1][30] ) );
  FDN1QM1P \Queue_reg[0][30]  ( .D(n475), .CPN(Clk_r), .Q(Packet_Out[30]) );
  FDN1QM1P \Queue_reg[1][29]  ( .D(n442), .CPN(Clk_r), .Q(\Queue[1][29] ) );
  FDN1QM1P \Queue_reg[0][29]  ( .D(n474), .CPN(Clk_r), .Q(Packet_Out[29]) );
  FDN1QM1P \Queue_reg[1][28]  ( .D(n441), .CPN(Clk_r), .Q(\Queue[1][28] ) );
  FDN1QM1P \Queue_reg[0][28]  ( .D(n473), .CPN(Clk_r), .Q(Packet_Out[28]) );
  FDN1QM1P \Queue_reg[1][27]  ( .D(n440), .CPN(Clk_r), .Q(\Queue[1][27] ) );
  FDN1QM1P \Queue_reg[0][27]  ( .D(n472), .CPN(Clk_r), .Q(Packet_Out[27]) );
  FDN1QM1P \Queue_reg[1][26]  ( .D(n439), .CPN(Clk_r), .Q(\Queue[1][26] ) );
  FDN1QM1P \Queue_reg[0][26]  ( .D(n471), .CPN(Clk_r), .Q(Packet_Out[26]) );
  FDN1QM1P \Queue_reg[1][25]  ( .D(n438), .CPN(Clk_r), .Q(\Queue[1][25] ) );
  FDN1QM1P \Queue_reg[0][25]  ( .D(n470), .CPN(Clk_r), .Q(Packet_Out[25]) );
  FDN1QM1P \Queue_reg[1][24]  ( .D(n437), .CPN(Clk_r), .Q(\Queue[1][24] ) );
  FDN1QM1P \Queue_reg[0][24]  ( .D(n469), .CPN(Clk_r), .Q(Packet_Out[24]) );
  FDN1QM1P \Queue_reg[1][23]  ( .D(n436), .CPN(Clk_r), .Q(\Queue[1][23] ) );
  FDN1QM1P \Queue_reg[0][23]  ( .D(n468), .CPN(Clk_r), .Q(Packet_Out[23]) );
  FDN1QM1P \Queue_reg[1][22]  ( .D(n435), .CPN(Clk_r), .Q(\Queue[1][22] ) );
  FDN1QM1P \Queue_reg[0][22]  ( .D(n467), .CPN(Clk_r), .Q(Packet_Out[22]) );
  FDN1QM1P \Queue_reg[1][21]  ( .D(n434), .CPN(Clk_r), .Q(\Queue[1][21] ) );
  FDN1QM1P \Queue_reg[0][21]  ( .D(n466), .CPN(Clk_r), .Q(Packet_Out[21]) );
  FDN1QM1P \Queue_reg[1][20]  ( .D(n433), .CPN(Clk_r), .Q(\Queue[1][20] ) );
  FDN1QM1P \Queue_reg[0][20]  ( .D(n465), .CPN(Clk_r), .Q(Packet_Out[20]) );
  FDN1QM1P \Queue_reg[1][19]  ( .D(n432), .CPN(Clk_r), .Q(\Queue[1][19] ) );
  FDN1QM1P \Queue_reg[0][19]  ( .D(n464), .CPN(Clk_r), .Q(Packet_Out[19]) );
  FDN1QM1P \Queue_reg[1][18]  ( .D(n431), .CPN(Clk_r), .Q(\Queue[1][18] ) );
  FDN1QM1P \Queue_reg[0][18]  ( .D(n463), .CPN(Clk_r), .Q(Packet_Out[18]) );
  FDN1QM1P \Queue_reg[1][17]  ( .D(n430), .CPN(Clk_r), .Q(\Queue[1][17] ) );
  FDN1QM1P \Queue_reg[0][17]  ( .D(n462), .CPN(Clk_r), .Q(Packet_Out[17]) );
  FDN1QM1P \Queue_reg[1][16]  ( .D(n429), .CPN(Clk_r), .Q(\Queue[1][16] ) );
  FDN1QM1P \Queue_reg[0][16]  ( .D(n461), .CPN(Clk_r), .Q(Packet_Out[16]) );
  FDN1QM1P \Queue_reg[1][15]  ( .D(n428), .CPN(Clk_r), .Q(\Queue[1][15] ) );
  FDN1QM1P \Queue_reg[0][15]  ( .D(n460), .CPN(Clk_r), .Q(Packet_Out[15]) );
  FDN1QM1P \Queue_reg[1][14]  ( .D(n427), .CPN(Clk_r), .Q(\Queue[1][14] ) );
  FDN1QM1P \Queue_reg[0][14]  ( .D(n459), .CPN(Clk_r), .Q(Packet_Out[14]) );
  FDN1QM1P \Queue_reg[1][13]  ( .D(n426), .CPN(Clk_r), .Q(\Queue[1][13] ) );
  FDN1QM1P \Queue_reg[0][13]  ( .D(n458), .CPN(Clk_r), .Q(Packet_Out[13]) );
  FDN1QM1P \Queue_reg[1][12]  ( .D(n425), .CPN(Clk_r), .Q(\Queue[1][12] ) );
  FDN1QM1P \Queue_reg[0][12]  ( .D(n457), .CPN(Clk_r), .Q(Packet_Out[12]) );
  FDN1QM1P \Queue_reg[1][11]  ( .D(n424), .CPN(Clk_r), .Q(\Queue[1][11] ) );
  FDN1QM1P \Queue_reg[0][11]  ( .D(n456), .CPN(Clk_r), .Q(Packet_Out[11]) );
  FDN1QM1P \Queue_reg[1][10]  ( .D(n423), .CPN(Clk_r), .Q(\Queue[1][10] ) );
  FDN1QM1P \Queue_reg[0][10]  ( .D(n455), .CPN(Clk_r), .Q(Packet_Out[10]) );
  FDN1QM1P \Queue_reg[1][9]  ( .D(n422), .CPN(Clk_r), .Q(\Queue[1][9] ) );
  FDN1QM1P \Queue_reg[0][9]  ( .D(n454), .CPN(Clk_r), .Q(Packet_Out[9]) );
  FDN1QM1P \Queue_reg[1][8]  ( .D(n421), .CPN(Clk_r), .Q(\Queue[1][8] ) );
  FDN1QM1P \Queue_reg[0][8]  ( .D(n453), .CPN(Clk_r), .Q(Packet_Out[8]) );
  FDN1QM1P \Queue_reg[1][7]  ( .D(n420), .CPN(Clk_r), .Q(\Queue[1][7] ) );
  FDN1QM1P \Queue_reg[0][7]  ( .D(n452), .CPN(Clk_r), .Q(Packet_Out[7]) );
  FDN1QM1P \Queue_reg[1][6]  ( .D(n419), .CPN(Clk_r), .Q(\Queue[1][6] ) );
  FDN1QM1P \Queue_reg[0][6]  ( .D(n451), .CPN(Clk_r), .Q(Packet_Out[6]) );
  FDN1QM1P \Queue_reg[1][5]  ( .D(n418), .CPN(Clk_r), .Q(\Queue[1][5] ) );
  FDN1QM1P \Queue_reg[0][5]  ( .D(n450), .CPN(Clk_r), .Q(Packet_Out[5]) );
  FDN1QM1P \Queue_reg[1][4]  ( .D(n417), .CPN(Clk_r), .Q(\Queue[1][4] ) );
  FDN1QM1P \Queue_reg[0][4]  ( .D(n449), .CPN(Clk_r), .Q(Packet_Out[4]) );
  FDN1QM1P \Queue_reg[1][3]  ( .D(n416), .CPN(Clk_r), .Q(\Queue[1][3] ) );
  FDN1QM1P \Queue_reg[0][3]  ( .D(n448), .CPN(Clk_r), .Q(Packet_Out[3]) );
  FDN1QM1P \Queue_reg[1][2]  ( .D(n415), .CPN(Clk_r), .Q(\Queue[1][2] ) );
  FDN1QM1P \Queue_reg[0][2]  ( .D(n447), .CPN(Clk_r), .Q(Packet_Out[2]) );
  FDN1QM1P \Queue_reg[1][1]  ( .D(n414), .CPN(Clk_r), .Q(\Queue[1][1] ) );
  FDN1QM1P \Queue_reg[0][1]  ( .D(n446), .CPN(Clk_r), .Q(Packet_Out[1]) );
  FDN1QM1P \Queue_reg[1][0]  ( .D(n413), .CPN(Clk_r), .Q(\Queue[1][0] ) );
  FDN1QM1P \Queue_reg[0][0]  ( .D(n445), .CPN(Clk_r), .Q(Packet_Out[0]) );
  FDN2QM1P Empty_reg ( .D(n542), .CPN(Clk_r), .CD(Rst_n), .Q(n541) );
  NR3M1P U3 ( .A(Count[0]), .B(Count[2]), .C(n22), .Z(n100) );
  BUFM2P U4 ( .A(n97), .Z(n9) );
  BUFM1P U5 ( .A(n97), .Z(n10) );
  BUFM1P U6 ( .A(n205), .Z(n12) );
  BUFM2P U7 ( .A(n132), .Z(n3) );
  BUFM1P U8 ( .A(n205), .Z(n11) );
  NR2FM1P U9 ( .A(Read_Ack), .B(n99), .Z(n18) );
  NR3M1P U10 ( .A(n23), .B(Count[2]), .C(Count[1]), .Z(n376) );
  N1M1P U11 ( .A(Read_Ack), .Z(n137) );
  NR3M1P U12 ( .A(Count[2]), .B(n23), .C(n22), .Z(n140) );
  AOI21M2P U13 ( .A(n4), .B(n376), .C(n141), .Z(n95) );
  AOI21M3P U14 ( .A(n4), .B(n100), .C(n141), .Z(n57) );
  OAI211M4P U15 ( .A(n100), .B(n137), .C(n4), .D(n24), .Z(n59) );
  NR2FM3P U16 ( .A(n61), .B(n21), .Z(n20) );
  OAI211M4P U17 ( .A(n142), .B(n137), .C(n4), .D(n136), .Z(n208) );
  OAI211M4P U18 ( .A(n140), .B(n137), .C(n4), .D(n98), .Z(n135) );
  OAI21M2P U19 ( .A(n4), .B(Read_Ack), .C(n24), .Z(n56) );
  N1M2P U20 ( .A(n4), .Z(n99) );
  N1M1P U21 ( .A(n142), .Z(n21) );
  NR3M1P U22 ( .A(Count[0]), .B(Count[1]), .C(n19), .Z(n142) );
  N1M1P U23 ( .A(Count[1]), .Z(n22) );
  N1M1P U24 ( .A(Count[2]), .Z(n19) );
  N1M1P U25 ( .A(Count[0]), .Z(n23) );
  BUFM2P U26 ( .A(n95), .Z(n8) );
  AOI21M6P U27 ( .A(n4), .B(n142), .C(n141), .Z(n205) );
  ND2M2P U28 ( .A(Read_Ack), .B(Rst_n), .Z(n141) );
  ND2M2P U29 ( .A(n18), .B(Rst_n), .Z(n61) );
  BUFM10P U30 ( .A(Write_Ack), .Z(n4) );
  OAI211M4P U31 ( .A(n100), .B(n139), .C(Rst_n), .D(n138), .Z(n133) );
  N1M1P U32 ( .A(Packet_In[31]), .Z(n373) );
  N1M1P U33 ( .A(Packet_In[23]), .Z(n190) );
  N1M1P U34 ( .A(Packet_In[28]), .Z(n200) );
  N1M1P U35 ( .A(Packet_In[25]), .Z(n194) );
  N1M1P U36 ( .A(Packet_In[27]), .Z(n198) );
  N1M1P U37 ( .A(Packet_In[29]), .Z(n202) );
  N1M1P U38 ( .A(Packet_In[26]), .Z(n196) );
  OAI211M4P U39 ( .A(n140), .B(n139), .C(Rst_n), .D(n138), .Z(n206) );
  N1M1P U40 ( .A(Packet_In[24]), .Z(n192) );
  N1M1P U41 ( .A(Packet_In[21]), .Z(n186) );
  N1M1P U42 ( .A(Packet_In[22]), .Z(n188) );
  N1M1P U43 ( .A(Packet_In[20]), .Z(n184) );
  N1M1P U44 ( .A(Packet_In[19]), .Z(n182) );
  N1M1P U45 ( .A(Packet_In[7]), .Z(n158) );
  N1M1P U46 ( .A(Packet_In[8]), .Z(n160) );
  N1M1P U47 ( .A(Packet_In[30]), .Z(n204) );
  N1M1P U48 ( .A(Packet_In[2]), .Z(n148) );
  N1M1P U49 ( .A(Packet_In[5]), .Z(n154) );
  N1M1P U50 ( .A(Packet_In[14]), .Z(n172) );
  N1M1P U51 ( .A(Packet_In[16]), .Z(n176) );
  N1M1P U52 ( .A(Packet_In[0]), .Z(n144) );
  N1M1P U53 ( .A(Packet_In[6]), .Z(n156) );
  N1M1P U54 ( .A(Packet_In[4]), .Z(n152) );
  N1M1P U55 ( .A(Packet_In[15]), .Z(n174) );
  N1M1P U56 ( .A(Packet_In[18]), .Z(n180) );
  N1M1P U57 ( .A(Packet_In[12]), .Z(n168) );
  N1M1P U58 ( .A(Packet_In[1]), .Z(n146) );
  N1M1P U59 ( .A(Packet_In[3]), .Z(n150) );
  N1M1P U60 ( .A(Packet_In[11]), .Z(n166) );
  N1M1P U61 ( .A(Packet_In[10]), .Z(n164) );
  N1M1P U62 ( .A(Packet_In[17]), .Z(n178) );
  N1M1P U63 ( .A(Packet_In[13]), .Z(n170) );
  N1M1P U64 ( .A(Packet_In[9]), .Z(n162) );
  BUFM2P U65 ( .A(n57), .Z(n7) );
  BUFM2P U66 ( .A(n56), .Z(n6) );
  BUFM2P U67 ( .A(n56), .Z(n5) );
  N1M2P U68 ( .A(n18), .Z(n139) );
  N1M2P U69 ( .A(n62), .Z(n94) );
  OAI211M1P U70 ( .A(n376), .B(n137), .C(n4), .D(n62), .Z(n97) );
  NR2M1P U71 ( .A(n137), .B(n4), .Z(n375) );
  NR2M1P U72 ( .A(n18), .B(n375), .Z(n374) );
  AOI22CDNM1P U73 ( .A(n374), .B(n23), .C(n374), .D(n23), .Z(n377) );
  N1M1P U74 ( .A(n375), .Z(n17) );
  AOI22M1P U75 ( .A(Count[0]), .B(n139), .C(n17), .D(n23), .Z(n14) );
  AOI22CDNM1P U76 ( .A(Count[1]), .B(n14), .C(n14), .D(Count[1]), .Z(n378) );
  ND3M1P U77 ( .A(n23), .B(n19), .C(n22), .Z(n60) );
  ND2M1P U78 ( .A(Count[1]), .B(Read_Ack), .Z(n13) );
  OAI211M1P U79 ( .A(Count[1]), .B(n139), .C(n14), .D(n13), .Z(n15) );
  AOI22M1P U80 ( .A(n18), .B(n140), .C(Count[2]), .D(n15), .Z(n16) );
  OAI21M1P U81 ( .A(n60), .B(n17), .C(n16), .Z(n379) );
  AOI22CDNM1P U82 ( .A(n20), .B(n373), .C(\Queue[4][31] ), .D(n20), .Z(n380)
         );
  AOI22CDNM1P U83 ( .A(n20), .B(n144), .C(\Queue[4][0] ), .D(n20), .Z(n381) );
  AOI22CDNM1P U84 ( .A(n20), .B(n146), .C(\Queue[4][1] ), .D(n20), .Z(n382) );
  AOI22CDNM1P U85 ( .A(n20), .B(n148), .C(\Queue[4][2] ), .D(n20), .Z(n383) );
  AOI22CDNM1P U86 ( .A(n20), .B(n150), .C(\Queue[4][3] ), .D(n20), .Z(n384) );
  AOI22CDNM1P U87 ( .A(n20), .B(n152), .C(\Queue[4][4] ), .D(n20), .Z(n385) );
  AOI22CDNM1P U88 ( .A(n20), .B(n154), .C(\Queue[4][5] ), .D(n20), .Z(n386) );
  AOI22CDNM1P U89 ( .A(n20), .B(n156), .C(\Queue[4][6] ), .D(n20), .Z(n387) );
  AOI22CDNM1P U90 ( .A(n20), .B(n158), .C(\Queue[4][7] ), .D(n20), .Z(n388) );
  AOI22CDNM1P U91 ( .A(n20), .B(n160), .C(\Queue[4][8] ), .D(n20), .Z(n389) );
  AOI22CDNM1P U92 ( .A(n20), .B(n162), .C(\Queue[4][9] ), .D(n20), .Z(n390) );
  AOI22CDNM1P U93 ( .A(n20), .B(n164), .C(\Queue[4][10] ), .D(n20), .Z(n391)
         );
  AOI22CDNM1P U94 ( .A(n20), .B(n166), .C(\Queue[4][11] ), .D(n20), .Z(n392)
         );
  AOI22CDNM1P U95 ( .A(n20), .B(n168), .C(\Queue[4][12] ), .D(n20), .Z(n393)
         );
  AOI22CDNM1P U96 ( .A(n20), .B(n170), .C(\Queue[4][13] ), .D(n20), .Z(n394)
         );
  AOI22CDNM1P U97 ( .A(n20), .B(n172), .C(\Queue[4][14] ), .D(n20), .Z(n395)
         );
  AOI22CDNM1P U98 ( .A(n20), .B(n174), .C(\Queue[4][15] ), .D(n20), .Z(n396)
         );
  AOI22CDNM1P U99 ( .A(n20), .B(n176), .C(\Queue[4][16] ), .D(n20), .Z(n397)
         );
  AOI22CDNM1P U100 ( .A(n20), .B(n178), .C(\Queue[4][17] ), .D(n20), .Z(n398)
         );
  AOI22CDNM1P U101 ( .A(n20), .B(n180), .C(\Queue[4][18] ), .D(n20), .Z(n399)
         );
  AOI22CDNM1P U102 ( .A(n20), .B(n182), .C(\Queue[4][19] ), .D(n20), .Z(n400)
         );
  AOI22CDNM1P U103 ( .A(n20), .B(n184), .C(\Queue[4][20] ), .D(n20), .Z(n401)
         );
  AOI22CDNM1P U104 ( .A(n20), .B(n186), .C(\Queue[4][21] ), .D(n20), .Z(n402)
         );
  AOI22CDNM1P U105 ( .A(n20), .B(n188), .C(\Queue[4][22] ), .D(n20), .Z(n403)
         );
  AOI22CDNM1P U106 ( .A(n20), .B(n190), .C(\Queue[4][23] ), .D(n20), .Z(n404)
         );
  AOI22CDNM1P U107 ( .A(n20), .B(n192), .C(\Queue[4][24] ), .D(n20), .Z(n405)
         );
  AOI22CDNM1P U108 ( .A(n20), .B(n194), .C(\Queue[4][25] ), .D(n20), .Z(n406)
         );
  AOI22CDNM1P U109 ( .A(n20), .B(n196), .C(\Queue[4][26] ), .D(n20), .Z(n407)
         );
  AOI22CDNM1P U110 ( .A(n20), .B(n198), .C(\Queue[4][27] ), .D(n20), .Z(n408)
         );
  AOI22CDNM1P U111 ( .A(n20), .B(n200), .C(\Queue[4][28] ), .D(n20), .Z(n409)
         );
  AOI22CDNM1P U112 ( .A(n20), .B(n202), .C(\Queue[4][29] ), .D(n20), .Z(n410)
         );
  AOI22CDNM1P U113 ( .A(n20), .B(n204), .C(\Queue[4][30] ), .D(n20), .Z(n411)
         );
  OAI22CDNM1P U114 ( .A(n139), .B(n21), .C(n374), .D(Full), .Z(n412) );
  OA21M1P U115 ( .A(n139), .B(n376), .C(Rst_n), .Z(n24) );
  AOI22M1P U116 ( .A(\Queue[2][0] ), .B(n57), .C(\Queue[1][0] ), .D(n5), .Z(
        n25) );
  OAI21M1P U117 ( .A(n144), .B(n59), .C(n25), .Z(n413) );
  AOI22M1P U118 ( .A(n7), .B(\Queue[2][1] ), .C(\Queue[1][1] ), .D(n5), .Z(n26) );
  OAI21M1P U119 ( .A(n59), .B(n146), .C(n26), .Z(n414) );
  AOI22M1P U120 ( .A(n57), .B(\Queue[2][2] ), .C(\Queue[1][2] ), .D(n5), .Z(
        n27) );
  OAI21M1P U121 ( .A(n59), .B(n148), .C(n27), .Z(n415) );
  AOI22M1P U122 ( .A(n57), .B(\Queue[2][3] ), .C(\Queue[1][3] ), .D(n5), .Z(
        n28) );
  OAI21M1P U123 ( .A(n59), .B(n150), .C(n28), .Z(n416) );
  AOI22M1P U124 ( .A(n57), .B(\Queue[2][4] ), .C(\Queue[1][4] ), .D(n5), .Z(
        n29) );
  OAI21M1P U125 ( .A(n59), .B(n152), .C(n29), .Z(n417) );
  AOI22M1P U126 ( .A(n57), .B(\Queue[2][5] ), .C(\Queue[1][5] ), .D(n5), .Z(
        n30) );
  OAI21M1P U127 ( .A(n59), .B(n154), .C(n30), .Z(n418) );
  AOI22M1P U128 ( .A(n57), .B(\Queue[2][6] ), .C(\Queue[1][6] ), .D(n5), .Z(
        n31) );
  OAI21M1P U129 ( .A(n59), .B(n156), .C(n31), .Z(n419) );
  AOI22M1P U130 ( .A(n57), .B(\Queue[2][7] ), .C(\Queue[1][7] ), .D(n5), .Z(
        n32) );
  OAI21M1P U131 ( .A(n59), .B(n158), .C(n32), .Z(n420) );
  AOI22M1P U132 ( .A(n57), .B(\Queue[2][8] ), .C(\Queue[1][8] ), .D(n5), .Z(
        n33) );
  OAI21M1P U133 ( .A(n59), .B(n160), .C(n33), .Z(n421) );
  AOI22M1P U134 ( .A(n7), .B(\Queue[2][9] ), .C(\Queue[1][9] ), .D(n56), .Z(
        n34) );
  OAI21M1P U135 ( .A(n59), .B(n162), .C(n34), .Z(n422) );
  AOI22M1P U136 ( .A(n57), .B(\Queue[2][10] ), .C(\Queue[1][10] ), .D(n5), .Z(
        n35) );
  OAI21M1P U137 ( .A(n59), .B(n164), .C(n35), .Z(n423) );
  AOI22M1P U138 ( .A(n57), .B(\Queue[2][11] ), .C(\Queue[1][11] ), .D(n6), .Z(
        n36) );
  OAI21M1P U139 ( .A(n59), .B(n166), .C(n36), .Z(n424) );
  AOI22M1P U140 ( .A(n7), .B(\Queue[2][12] ), .C(\Queue[1][12] ), .D(n56), .Z(
        n37) );
  OAI21M1P U141 ( .A(n59), .B(n168), .C(n37), .Z(n425) );
  AOI22M1P U142 ( .A(n7), .B(\Queue[2][13] ), .C(\Queue[1][13] ), .D(n56), .Z(
        n38) );
  OAI21M1P U143 ( .A(n59), .B(n170), .C(n38), .Z(n426) );
  AOI22M1P U144 ( .A(n7), .B(\Queue[2][14] ), .C(\Queue[1][14] ), .D(n56), .Z(
        n39) );
  OAI21M1P U145 ( .A(n59), .B(n172), .C(n39), .Z(n427) );
  AOI22M1P U146 ( .A(n7), .B(\Queue[2][15] ), .C(\Queue[1][15] ), .D(n56), .Z(
        n40) );
  OAI21M1P U147 ( .A(n59), .B(n174), .C(n40), .Z(n428) );
  AOI22M1P U148 ( .A(n7), .B(\Queue[2][16] ), .C(\Queue[1][16] ), .D(n56), .Z(
        n41) );
  OAI21M1P U149 ( .A(n59), .B(n176), .C(n41), .Z(n429) );
  AOI22M1P U150 ( .A(n7), .B(\Queue[2][17] ), .C(\Queue[1][17] ), .D(n56), .Z(
        n42) );
  OAI21M1P U151 ( .A(n59), .B(n178), .C(n42), .Z(n430) );
  AOI22M1P U152 ( .A(n7), .B(\Queue[2][18] ), .C(\Queue[1][18] ), .D(n6), .Z(
        n43) );
  OAI21M1P U153 ( .A(n59), .B(n180), .C(n43), .Z(n431) );
  AOI22M1P U154 ( .A(n7), .B(\Queue[2][19] ), .C(\Queue[1][19] ), .D(n6), .Z(
        n44) );
  OAI21M1P U155 ( .A(n59), .B(n182), .C(n44), .Z(n432) );
  AOI22M1P U156 ( .A(n7), .B(\Queue[2][20] ), .C(\Queue[1][20] ), .D(n6), .Z(
        n45) );
  OAI21M1P U157 ( .A(n59), .B(n184), .C(n45), .Z(n433) );
  AOI22M1P U158 ( .A(n7), .B(\Queue[2][21] ), .C(\Queue[1][21] ), .D(n6), .Z(
        n46) );
  OAI21M1P U159 ( .A(n59), .B(n186), .C(n46), .Z(n434) );
  AOI22M1P U160 ( .A(n57), .B(\Queue[2][22] ), .C(\Queue[1][22] ), .D(n6), .Z(
        n47) );
  OAI21M1P U161 ( .A(n59), .B(n188), .C(n47), .Z(n435) );
  AOI22M1P U162 ( .A(n7), .B(\Queue[2][23] ), .C(\Queue[1][23] ), .D(n6), .Z(
        n48) );
  OAI21M1P U163 ( .A(n59), .B(n190), .C(n48), .Z(n436) );
  AOI22M1P U164 ( .A(n57), .B(\Queue[2][24] ), .C(\Queue[1][24] ), .D(n6), .Z(
        n49) );
  OAI21M1P U165 ( .A(n59), .B(n192), .C(n49), .Z(n437) );
  AOI22M1P U166 ( .A(n57), .B(\Queue[2][25] ), .C(\Queue[1][25] ), .D(n6), .Z(
        n50) );
  OAI21M1P U167 ( .A(n59), .B(n194), .C(n50), .Z(n438) );
  AOI22M1P U168 ( .A(n57), .B(\Queue[2][26] ), .C(\Queue[1][26] ), .D(n6), .Z(
        n51) );
  OAI21M1P U169 ( .A(n59), .B(n196), .C(n51), .Z(n439) );
  AOI22M1P U170 ( .A(n57), .B(\Queue[2][27] ), .C(\Queue[1][27] ), .D(n6), .Z(
        n52) );
  OAI21M1P U171 ( .A(n59), .B(n198), .C(n52), .Z(n440) );
  AOI22M1P U172 ( .A(n57), .B(\Queue[2][28] ), .C(\Queue[1][28] ), .D(n5), .Z(
        n53) );
  OAI21M1P U173 ( .A(n59), .B(n200), .C(n53), .Z(n441) );
  AOI22M1P U174 ( .A(n57), .B(\Queue[2][29] ), .C(\Queue[1][29] ), .D(n5), .Z(
        n54) );
  OAI21M1P U175 ( .A(n59), .B(n202), .C(n54), .Z(n442) );
  AOI22M1P U176 ( .A(n57), .B(\Queue[2][30] ), .C(\Queue[1][30] ), .D(n6), .Z(
        n55) );
  OAI21M1P U177 ( .A(n59), .B(n204), .C(n55), .Z(n443) );
  AOI22M1P U178 ( .A(n57), .B(\Queue[2][31] ), .C(\Queue[1][31] ), .D(n5), .Z(
        n58) );
  OAI21M1P U179 ( .A(n59), .B(n373), .C(n58), .Z(n444) );
  OAI21M1P U180 ( .A(n61), .B(n60), .C(n141), .Z(n62) );
  AOI22M1P U181 ( .A(\Queue[1][0] ), .B(n8), .C(n94), .D(Packet_Out[0]), .Z(
        n63) );
  OAI21M1P U182 ( .A(n144), .B(n9), .C(n63), .Z(n445) );
  AOI22M1P U183 ( .A(\Queue[1][1] ), .B(n8), .C(n94), .D(Packet_Out[1]), .Z(
        n64) );
  OAI21M1P U184 ( .A(n146), .B(n9), .C(n64), .Z(n446) );
  AOI22M1P U185 ( .A(\Queue[1][2] ), .B(n8), .C(n94), .D(Packet_Out[2]), .Z(
        n65) );
  OAI21M1P U186 ( .A(n148), .B(n9), .C(n65), .Z(n447) );
  AOI22M1P U187 ( .A(\Queue[1][3] ), .B(n95), .C(n94), .D(Packet_Out[3]), .Z(
        n66) );
  OAI21M1P U188 ( .A(n150), .B(n9), .C(n66), .Z(n448) );
  AOI22M1P U189 ( .A(\Queue[1][4] ), .B(n95), .C(n94), .D(Packet_Out[4]), .Z(
        n67) );
  OAI21M1P U190 ( .A(n152), .B(n9), .C(n67), .Z(n449) );
  AOI22M1P U191 ( .A(\Queue[1][5] ), .B(n95), .C(n94), .D(Packet_Out[5]), .Z(
        n68) );
  OAI21M1P U192 ( .A(n154), .B(n9), .C(n68), .Z(n450) );
  AOI22M1P U193 ( .A(\Queue[1][6] ), .B(n95), .C(n94), .D(Packet_Out[6]), .Z(
        n69) );
  OAI21M1P U194 ( .A(n156), .B(n9), .C(n69), .Z(n451) );
  AOI22M1P U195 ( .A(\Queue[1][7] ), .B(n95), .C(n94), .D(Packet_Out[7]), .Z(
        n70) );
  OAI21M1P U196 ( .A(n158), .B(n9), .C(n70), .Z(n452) );
  AOI22M1P U197 ( .A(\Queue[1][8] ), .B(n95), .C(n94), .D(Packet_Out[8]), .Z(
        n71) );
  OAI21M1P U198 ( .A(n160), .B(n9), .C(n71), .Z(n453) );
  AOI22M1P U199 ( .A(\Queue[1][9] ), .B(n95), .C(n94), .D(Packet_Out[9]), .Z(
        n72) );
  OAI21M1P U200 ( .A(n162), .B(n9), .C(n72), .Z(n454) );
  AOI22M1P U201 ( .A(\Queue[1][10] ), .B(n8), .C(n94), .D(Packet_Out[10]), .Z(
        n73) );
  OAI21M1P U202 ( .A(n164), .B(n9), .C(n73), .Z(n455) );
  AOI22M1P U203 ( .A(\Queue[1][11] ), .B(n8), .C(n94), .D(Packet_Out[11]), .Z(
        n74) );
  OAI21M1P U204 ( .A(n166), .B(n9), .C(n74), .Z(n456) );
  AOI22M1P U205 ( .A(\Queue[1][12] ), .B(n8), .C(n94), .D(Packet_Out[12]), .Z(
        n75) );
  OAI21M1P U206 ( .A(n168), .B(n9), .C(n75), .Z(n457) );
  AOI22M1P U207 ( .A(\Queue[1][13] ), .B(n8), .C(n94), .D(Packet_Out[13]), .Z(
        n76) );
  OAI21M1P U208 ( .A(n170), .B(n9), .C(n76), .Z(n458) );
  AOI22M1P U209 ( .A(\Queue[1][14] ), .B(n8), .C(n94), .D(Packet_Out[14]), .Z(
        n77) );
  OAI21M1P U210 ( .A(n172), .B(n9), .C(n77), .Z(n459) );
  AOI22M1P U211 ( .A(\Queue[1][15] ), .B(n8), .C(n94), .D(Packet_Out[15]), .Z(
        n78) );
  OAI21M1P U212 ( .A(n174), .B(n9), .C(n78), .Z(n460) );
  AOI22M1P U213 ( .A(\Queue[1][16] ), .B(n95), .C(n94), .D(Packet_Out[16]), 
        .Z(n79) );
  OAI21M1P U214 ( .A(n176), .B(n9), .C(n79), .Z(n461) );
  AOI22M1P U215 ( .A(\Queue[1][17] ), .B(n95), .C(n94), .D(Packet_Out[17]), 
        .Z(n80) );
  OAI21M1P U216 ( .A(n178), .B(n9), .C(n80), .Z(n462) );
  AOI22M1P U217 ( .A(\Queue[1][18] ), .B(n95), .C(n94), .D(Packet_Out[18]), 
        .Z(n81) );
  OAI21M1P U218 ( .A(n180), .B(n9), .C(n81), .Z(n463) );
  AOI22M1P U219 ( .A(\Queue[1][19] ), .B(n95), .C(n94), .D(Packet_Out[19]), 
        .Z(n82) );
  OAI21M1P U220 ( .A(n182), .B(n9), .C(n82), .Z(n464) );
  AOI22M1P U221 ( .A(\Queue[1][20] ), .B(n8), .C(n94), .D(Packet_Out[20]), .Z(
        n83) );
  OAI21M1P U222 ( .A(n184), .B(n10), .C(n83), .Z(n465) );
  AOI22M1P U223 ( .A(\Queue[1][21] ), .B(n8), .C(n94), .D(Packet_Out[21]), .Z(
        n84) );
  OAI21M1P U224 ( .A(n186), .B(n10), .C(n84), .Z(n466) );
  AOI22M1P U225 ( .A(\Queue[1][22] ), .B(n8), .C(n94), .D(Packet_Out[22]), .Z(
        n85) );
  OAI21M1P U226 ( .A(n188), .B(n10), .C(n85), .Z(n467) );
  AOI22M1P U227 ( .A(\Queue[1][23] ), .B(n8), .C(n94), .D(Packet_Out[23]), .Z(
        n86) );
  OAI21M1P U228 ( .A(n190), .B(n10), .C(n86), .Z(n468) );
  AOI22M1P U229 ( .A(\Queue[1][24] ), .B(n8), .C(n94), .D(Packet_Out[24]), .Z(
        n87) );
  OAI21M1P U230 ( .A(n192), .B(n10), .C(n87), .Z(n469) );
  AOI22M1P U231 ( .A(\Queue[1][25] ), .B(n8), .C(n94), .D(Packet_Out[25]), .Z(
        n88) );
  OAI21M1P U232 ( .A(n194), .B(n10), .C(n88), .Z(n470) );
  AOI22M1P U233 ( .A(\Queue[1][26] ), .B(n8), .C(n94), .D(Packet_Out[26]), .Z(
        n89) );
  OAI21M1P U234 ( .A(n196), .B(n10), .C(n89), .Z(n471) );
  AOI22M1P U235 ( .A(\Queue[1][27] ), .B(n8), .C(n94), .D(Packet_Out[27]), .Z(
        n90) );
  OAI21M1P U236 ( .A(n198), .B(n10), .C(n90), .Z(n472) );
  AOI22M1P U237 ( .A(\Queue[1][28] ), .B(n8), .C(n94), .D(Packet_Out[28]), .Z(
        n91) );
  OAI21M1P U238 ( .A(n200), .B(n10), .C(n91), .Z(n473) );
  AOI22M1P U239 ( .A(\Queue[1][29] ), .B(n8), .C(n94), .D(Packet_Out[29]), .Z(
        n92) );
  OAI21M1P U240 ( .A(n202), .B(n10), .C(n92), .Z(n474) );
  AOI22M1P U241 ( .A(\Queue[1][30] ), .B(n95), .C(n94), .D(Packet_Out[30]), 
        .Z(n93) );
  OAI21M1P U242 ( .A(n204), .B(n9), .C(n93), .Z(n475) );
  AOI22M1P U243 ( .A(\Queue[1][31] ), .B(n8), .C(n94), .D(Packet_Out[31]), .Z(
        n96) );
  OAI21M1P U244 ( .A(n373), .B(n10), .C(n96), .Z(n476) );
  OA21M1P U245 ( .A(n139), .B(n100), .C(Rst_n), .Z(n98) );
  ND2M1P U246 ( .A(n99), .B(n137), .Z(n138) );
  AOI21M1P U247 ( .A(n4), .B(n140), .C(n141), .Z(n132) );
  AOI22M1P U248 ( .A(\Queue[2][0] ), .B(n133), .C(\Queue[3][0] ), .D(n3), .Z(
        n101) );
  OAI21M1P U249 ( .A(n144), .B(n135), .C(n101), .Z(n477) );
  AOI22M1P U250 ( .A(\Queue[2][1] ), .B(n133), .C(n3), .D(\Queue[3][1] ), .Z(
        n102) );
  OAI21M1P U251 ( .A(n146), .B(n135), .C(n102), .Z(n478) );
  AOI22M1P U252 ( .A(\Queue[2][2] ), .B(n133), .C(n3), .D(\Queue[3][2] ), .Z(
        n103) );
  OAI21M1P U253 ( .A(n148), .B(n135), .C(n103), .Z(n479) );
  AOI22M1P U254 ( .A(\Queue[2][3] ), .B(n133), .C(n3), .D(\Queue[3][3] ), .Z(
        n104) );
  OAI21M1P U255 ( .A(n150), .B(n135), .C(n104), .Z(n480) );
  AOI22M1P U256 ( .A(\Queue[2][4] ), .B(n133), .C(n3), .D(\Queue[3][4] ), .Z(
        n105) );
  OAI21M1P U257 ( .A(n152), .B(n135), .C(n105), .Z(n481) );
  AOI22M1P U258 ( .A(\Queue[2][5] ), .B(n133), .C(n3), .D(\Queue[3][5] ), .Z(
        n106) );
  OAI21M1P U259 ( .A(n154), .B(n135), .C(n106), .Z(n482) );
  AOI22M1P U260 ( .A(\Queue[2][6] ), .B(n133), .C(n3), .D(\Queue[3][6] ), .Z(
        n107) );
  OAI21M1P U261 ( .A(n156), .B(n135), .C(n107), .Z(n483) );
  AOI22M1P U262 ( .A(\Queue[2][7] ), .B(n133), .C(n3), .D(\Queue[3][7] ), .Z(
        n108) );
  OAI21M1P U263 ( .A(n158), .B(n135), .C(n108), .Z(n484) );
  AOI22M1P U264 ( .A(\Queue[2][8] ), .B(n133), .C(n3), .D(\Queue[3][8] ), .Z(
        n109) );
  OAI21M1P U265 ( .A(n160), .B(n135), .C(n109), .Z(n485) );
  AOI22M1P U266 ( .A(\Queue[2][9] ), .B(n133), .C(n3), .D(\Queue[3][9] ), .Z(
        n110) );
  OAI21M1P U267 ( .A(n162), .B(n135), .C(n110), .Z(n486) );
  AOI22M1P U268 ( .A(\Queue[2][10] ), .B(n133), .C(n3), .D(\Queue[3][10] ), 
        .Z(n111) );
  OAI21M1P U269 ( .A(n164), .B(n135), .C(n111), .Z(n487) );
  AOI22M1P U270 ( .A(\Queue[2][11] ), .B(n133), .C(n3), .D(\Queue[3][11] ), 
        .Z(n112) );
  OAI21M1P U271 ( .A(n166), .B(n135), .C(n112), .Z(n488) );
  AOI22M1P U272 ( .A(\Queue[2][12] ), .B(n133), .C(n3), .D(\Queue[3][12] ), 
        .Z(n113) );
  OAI21M1P U273 ( .A(n168), .B(n135), .C(n113), .Z(n489) );
  AOI22M1P U274 ( .A(\Queue[2][13] ), .B(n133), .C(n3), .D(\Queue[3][13] ), 
        .Z(n114) );
  OAI21M1P U275 ( .A(n170), .B(n135), .C(n114), .Z(n490) );
  AOI22M1P U276 ( .A(\Queue[2][14] ), .B(n133), .C(n3), .D(\Queue[3][14] ), 
        .Z(n115) );
  OAI21M1P U277 ( .A(n172), .B(n135), .C(n115), .Z(n491) );
  AOI22M1P U278 ( .A(\Queue[2][15] ), .B(n133), .C(n3), .D(\Queue[3][15] ), 
        .Z(n116) );
  OAI21M1P U279 ( .A(n174), .B(n135), .C(n116), .Z(n492) );
  AOI22M1P U280 ( .A(\Queue[2][16] ), .B(n133), .C(n3), .D(\Queue[3][16] ), 
        .Z(n117) );
  OAI21M1P U281 ( .A(n176), .B(n135), .C(n117), .Z(n493) );
  AOI22M1P U282 ( .A(\Queue[2][17] ), .B(n133), .C(n3), .D(\Queue[3][17] ), 
        .Z(n118) );
  OAI21M1P U283 ( .A(n178), .B(n135), .C(n118), .Z(n494) );
  AOI22M1P U284 ( .A(\Queue[2][18] ), .B(n133), .C(n3), .D(\Queue[3][18] ), 
        .Z(n119) );
  OAI21M1P U285 ( .A(n180), .B(n135), .C(n119), .Z(n495) );
  AOI22M1P U286 ( .A(\Queue[2][19] ), .B(n133), .C(n3), .D(\Queue[3][19] ), 
        .Z(n120) );
  OAI21M1P U287 ( .A(n182), .B(n135), .C(n120), .Z(n496) );
  AOI22M1P U288 ( .A(\Queue[2][20] ), .B(n133), .C(n3), .D(\Queue[3][20] ), 
        .Z(n121) );
  OAI21M1P U289 ( .A(n184), .B(n135), .C(n121), .Z(n497) );
  AOI22M1P U290 ( .A(\Queue[2][21] ), .B(n133), .C(n3), .D(\Queue[3][21] ), 
        .Z(n122) );
  OAI21M1P U291 ( .A(n186), .B(n135), .C(n122), .Z(n498) );
  AOI22M1P U292 ( .A(\Queue[2][22] ), .B(n133), .C(n3), .D(\Queue[3][22] ), 
        .Z(n123) );
  OAI21M1P U293 ( .A(n188), .B(n135), .C(n123), .Z(n499) );
  AOI22M1P U294 ( .A(\Queue[2][23] ), .B(n133), .C(n3), .D(\Queue[3][23] ), 
        .Z(n124) );
  OAI21M1P U295 ( .A(n190), .B(n135), .C(n124), .Z(n500) );
  AOI22M1P U296 ( .A(\Queue[2][24] ), .B(n133), .C(n3), .D(\Queue[3][24] ), 
        .Z(n125) );
  OAI21M1P U297 ( .A(n192), .B(n135), .C(n125), .Z(n501) );
  AOI22M1P U298 ( .A(\Queue[2][25] ), .B(n133), .C(n3), .D(\Queue[3][25] ), 
        .Z(n126) );
  OAI21M1P U299 ( .A(n194), .B(n135), .C(n126), .Z(n502) );
  AOI22M1P U300 ( .A(\Queue[2][26] ), .B(n133), .C(n3), .D(\Queue[3][26] ), 
        .Z(n127) );
  OAI21M1P U301 ( .A(n196), .B(n135), .C(n127), .Z(n503) );
  AOI22M1P U302 ( .A(\Queue[2][27] ), .B(n133), .C(n3), .D(\Queue[3][27] ), 
        .Z(n128) );
  OAI21M1P U303 ( .A(n198), .B(n135), .C(n128), .Z(n504) );
  AOI22M1P U304 ( .A(\Queue[2][28] ), .B(n133), .C(n3), .D(\Queue[3][28] ), 
        .Z(n129) );
  OAI21M1P U305 ( .A(n200), .B(n135), .C(n129), .Z(n505) );
  AOI22M1P U306 ( .A(\Queue[2][29] ), .B(n133), .C(n3), .D(\Queue[3][29] ), 
        .Z(n130) );
  OAI21M1P U307 ( .A(n202), .B(n135), .C(n130), .Z(n506) );
  AOI22M1P U308 ( .A(\Queue[2][30] ), .B(n133), .C(n3), .D(\Queue[3][30] ), 
        .Z(n131) );
  OAI21M1P U309 ( .A(n204), .B(n135), .C(n131), .Z(n507) );
  AOI22M1P U310 ( .A(\Queue[2][31] ), .B(n133), .C(n3), .D(\Queue[3][31] ), 
        .Z(n134) );
  OAI21M1P U311 ( .A(n373), .B(n135), .C(n134), .Z(n508) );
  OA21M1P U312 ( .A(n139), .B(n140), .C(Rst_n), .Z(n136) );
  AOI22M1P U313 ( .A(\Queue[3][0] ), .B(n206), .C(n205), .D(\Queue[4][0] ), 
        .Z(n143) );
  OAI21M1P U314 ( .A(n144), .B(n208), .C(n143), .Z(n509) );
  AOI22M1P U315 ( .A(\Queue[3][1] ), .B(n206), .C(n205), .D(\Queue[4][1] ), 
        .Z(n145) );
  OAI21M1P U316 ( .A(n146), .B(n208), .C(n145), .Z(n510) );
  AOI22M1P U317 ( .A(\Queue[3][2] ), .B(n206), .C(n205), .D(\Queue[4][2] ), 
        .Z(n147) );
  OAI21M1P U318 ( .A(n148), .B(n208), .C(n147), .Z(n511) );
  AOI22M1P U319 ( .A(\Queue[3][3] ), .B(n206), .C(n205), .D(\Queue[4][3] ), 
        .Z(n149) );
  OAI21M1P U320 ( .A(n150), .B(n208), .C(n149), .Z(n512) );
  AOI22M1P U321 ( .A(\Queue[3][4] ), .B(n206), .C(n205), .D(\Queue[4][4] ), 
        .Z(n151) );
  OAI21M1P U322 ( .A(n152), .B(n208), .C(n151), .Z(n513) );
  AOI22M1P U323 ( .A(\Queue[3][5] ), .B(n206), .C(n205), .D(\Queue[4][5] ), 
        .Z(n153) );
  OAI21M1P U324 ( .A(n154), .B(n208), .C(n153), .Z(n514) );
  AOI22M1P U325 ( .A(\Queue[3][6] ), .B(n206), .C(n205), .D(\Queue[4][6] ), 
        .Z(n155) );
  OAI21M1P U326 ( .A(n156), .B(n208), .C(n155), .Z(n515) );
  AOI22M1P U327 ( .A(\Queue[3][7] ), .B(n206), .C(n205), .D(\Queue[4][7] ), 
        .Z(n157) );
  OAI21M1P U328 ( .A(n158), .B(n208), .C(n157), .Z(n516) );
  AOI22M1P U329 ( .A(\Queue[3][8] ), .B(n206), .C(n11), .D(\Queue[4][8] ), .Z(
        n159) );
  OAI21M1P U330 ( .A(n160), .B(n208), .C(n159), .Z(n517) );
  AOI22M1P U331 ( .A(\Queue[3][9] ), .B(n206), .C(n12), .D(\Queue[4][9] ), .Z(
        n161) );
  OAI21M1P U332 ( .A(n162), .B(n208), .C(n161), .Z(n518) );
  AOI22M1P U333 ( .A(\Queue[3][10] ), .B(n206), .C(n11), .D(\Queue[4][10] ), 
        .Z(n163) );
  OAI21M1P U334 ( .A(n164), .B(n208), .C(n163), .Z(n519) );
  AOI22M1P U335 ( .A(\Queue[3][11] ), .B(n206), .C(n11), .D(\Queue[4][11] ), 
        .Z(n165) );
  OAI21M1P U336 ( .A(n166), .B(n208), .C(n165), .Z(n520) );
  AOI22M1P U337 ( .A(\Queue[3][12] ), .B(n206), .C(n11), .D(\Queue[4][12] ), 
        .Z(n167) );
  OAI21M1P U338 ( .A(n168), .B(n208), .C(n167), .Z(n521) );
  AOI22M1P U339 ( .A(\Queue[3][13] ), .B(n206), .C(n11), .D(\Queue[4][13] ), 
        .Z(n169) );
  OAI21M1P U340 ( .A(n170), .B(n208), .C(n169), .Z(n522) );
  AOI22M1P U341 ( .A(\Queue[3][14] ), .B(n206), .C(n11), .D(\Queue[4][14] ), 
        .Z(n171) );
  OAI21M1P U342 ( .A(n172), .B(n208), .C(n171), .Z(n523) );
  AOI22M1P U343 ( .A(\Queue[3][15] ), .B(n206), .C(n11), .D(\Queue[4][15] ), 
        .Z(n173) );
  OAI21M1P U344 ( .A(n174), .B(n208), .C(n173), .Z(n524) );
  AOI22M1P U345 ( .A(\Queue[3][16] ), .B(n206), .C(n11), .D(\Queue[4][16] ), 
        .Z(n175) );
  OAI21M1P U346 ( .A(n176), .B(n208), .C(n175), .Z(n525) );
  AOI22M1P U347 ( .A(\Queue[3][17] ), .B(n206), .C(n11), .D(\Queue[4][17] ), 
        .Z(n177) );
  OAI21M1P U348 ( .A(n178), .B(n208), .C(n177), .Z(n526) );
  AOI22M1P U349 ( .A(\Queue[3][18] ), .B(n206), .C(n11), .D(\Queue[4][18] ), 
        .Z(n179) );
  OAI21M1P U350 ( .A(n180), .B(n208), .C(n179), .Z(n527) );
  AOI22M1P U351 ( .A(\Queue[3][19] ), .B(n206), .C(n11), .D(\Queue[4][19] ), 
        .Z(n181) );
  OAI21M1P U352 ( .A(n182), .B(n208), .C(n181), .Z(n528) );
  AOI22M1P U353 ( .A(\Queue[3][20] ), .B(n206), .C(n12), .D(\Queue[4][20] ), 
        .Z(n183) );
  OAI21M1P U354 ( .A(n184), .B(n208), .C(n183), .Z(n529) );
  AOI22M1P U355 ( .A(\Queue[3][21] ), .B(n206), .C(n12), .D(\Queue[4][21] ), 
        .Z(n185) );
  OAI21M1P U356 ( .A(n186), .B(n208), .C(n185), .Z(n530) );
  AOI22M1P U357 ( .A(\Queue[3][22] ), .B(n206), .C(n12), .D(\Queue[4][22] ), 
        .Z(n187) );
  OAI21M1P U358 ( .A(n188), .B(n208), .C(n187), .Z(n531) );
  AOI22M1P U359 ( .A(\Queue[3][23] ), .B(n206), .C(n12), .D(\Queue[4][23] ), 
        .Z(n189) );
  OAI21M1P U360 ( .A(n190), .B(n208), .C(n189), .Z(n532) );
  AOI22M1P U361 ( .A(\Queue[3][24] ), .B(n206), .C(n12), .D(\Queue[4][24] ), 
        .Z(n191) );
  OAI21M1P U362 ( .A(n192), .B(n208), .C(n191), .Z(n533) );
  AOI22M1P U363 ( .A(\Queue[3][25] ), .B(n206), .C(n12), .D(\Queue[4][25] ), 
        .Z(n193) );
  OAI21M1P U364 ( .A(n194), .B(n208), .C(n193), .Z(n534) );
  AOI22M1P U365 ( .A(\Queue[3][26] ), .B(n206), .C(n12), .D(\Queue[4][26] ), 
        .Z(n195) );
  OAI21M1P U366 ( .A(n196), .B(n208), .C(n195), .Z(n535) );
  AOI22M1P U367 ( .A(\Queue[3][27] ), .B(n206), .C(n12), .D(\Queue[4][27] ), 
        .Z(n197) );
  OAI21M1P U368 ( .A(n198), .B(n208), .C(n197), .Z(n536) );
  AOI22M1P U369 ( .A(\Queue[3][28] ), .B(n206), .C(n12), .D(\Queue[4][28] ), 
        .Z(n199) );
  OAI21M1P U370 ( .A(n200), .B(n208), .C(n199), .Z(n537) );
  AOI22M1P U371 ( .A(\Queue[3][29] ), .B(n206), .C(n12), .D(\Queue[4][29] ), 
        .Z(n201) );
  OAI21M1P U372 ( .A(n202), .B(n208), .C(n201), .Z(n538) );
  AOI22M1P U373 ( .A(\Queue[3][30] ), .B(n206), .C(n11), .D(\Queue[4][30] ), 
        .Z(n203) );
  OAI21M1P U374 ( .A(n204), .B(n208), .C(n203), .Z(n539) );
  AOI22M1P U375 ( .A(\Queue[3][31] ), .B(n206), .C(n12), .D(\Queue[4][31] ), 
        .Z(n207) );
  OAI21M1P U376 ( .A(n373), .B(n208), .C(n207), .Z(n540) );
  N1M1P U377 ( .A(n541), .Z(Empty) );
  AOI22M1P U378 ( .A(n376), .B(n375), .C(n374), .D(Empty), .Z(n542) );
endmodule


module Link_Control_3 ( Clk_r, Rst_n, Tx_Ready, Tx_Error, RxData_Valid, RxData, 
        Packet_From_Core, TxQueue_Write, RxQueue_Read, TxData_Valid, TxData, 
        Error_Ack, Core_Rcv_Ready, Packet_To_Core, RxQueue_Empty, TxQueue_Full
 );
  input [31:0] RxData;
  input [31:0] Packet_From_Core;
  output [31:0] TxData;
  output [31:0] Packet_To_Core;
  input Clk_r, Rst_n, Tx_Ready, Tx_Error, RxData_Valid, TxQueue_Write,
         RxQueue_Read;
  output TxData_Valid, Error_Ack, Core_Rcv_Ready, RxQueue_Empty, TxQueue_Full;
  wire   TxQueue_Read, TxQueue_Empty, RxQueue_Write, RxQueue_Full, N9, N16, n5,
         n6, n7, n8, n9;

  Packet_Queue_8 TxQueue ( .Clk_r(Clk_r), .Rst_n(Rst_n), .Packet_In(
        Packet_From_Core), .Read_Ack(TxQueue_Read), .Write_Ack(TxQueue_Write), 
        .Packet_Out(TxData), .Empty(TxQueue_Empty), .Full(TxQueue_Full) );
  Packet_Queue_7 RxQueue ( .Clk_r(Clk_r), .Rst_n(Rst_n), .Packet_In(RxData), 
        .Read_Ack(RxQueue_Read), .Write_Ack(RxQueue_Write), .Packet_Out(
        Packet_To_Core), .Empty(RxQueue_Empty), .Full(RxQueue_Full) );
  FD2QM1P Core_Rcv_Ready_reg ( .D(N9), .CP(Clk_r), .CD(Rst_n), .Q(
        Core_Rcv_Ready) );
  FD2QM1P TxQueue_Read_reg ( .D(N16), .CP(Clk_r), .CD(Rst_n), .Q(TxQueue_Read)
         );
  FD2QM1P Error_Ack_reg ( .D(Tx_Error), .CP(Clk_r), .CD(Rst_n), .Q(Error_Ack)
         );
  FD4QM1P RxQueue_Write_reg ( .D(n7), .CP(Clk_r), .SD(Rst_n), .Q(n6) );
  FD4QM1P TxData_Valid_reg ( .D(n9), .CP(Clk_r), .SD(Rst_n), .Q(n8) );
  N1M2P U3 ( .A(n6), .Z(RxQueue_Write) );
  NR2M1P U4 ( .A(n8), .B(Tx_Ready), .Z(N16) );
  NR2M1P U5 ( .A(RxData_Valid), .B(RxQueue_Full), .Z(n5) );
  OA21M1P U6 ( .A(Core_Rcv_Ready), .B(n5), .C(n6), .Z(N9) );
  N1M1P U7 ( .A(n8), .Z(TxData_Valid) );
  ND3M1P U8 ( .A(n6), .B(Core_Rcv_Ready), .C(RxData_Valid), .Z(n7) );
  AO21CNM1P U9 ( .A(n8), .B(TxQueue_Empty), .C(Tx_Ready), .Z(n9) );
endmodule


module core_synth ( Clk_r, Rst_n, N_Tx_Ready, N_Tx_Error, N_RxData_Valid, N_RxData, 
        S_Tx_Ready, S_Tx_Error, S_RxData_Valid, S_RxData, W_Tx_Ready, 
        W_Tx_Error, W_RxData_Valid, W_RxData, E_Tx_Ready, E_Tx_Error, 
        E_RxData_Valid, E_RxData, Packet_From_Node, Packet_From_Node_Valid, 
        N_TxData_Valid, N_TxData, N_Error_Ack, N_Core_Rcv_Ready, 
        S_TxData_Valid, S_TxData, S_Error_Ack, S_Core_Rcv_Ready, 
        W_TxData_Valid, W_TxData, W_Error_Ack, W_Core_Rcv_Ready, 
        E_TxData_Valid, E_TxData, E_Error_Ack, E_Core_Rcv_Ready, Core_Load_Ack, 
        Packet_To_Node, Packet_To_Node_Valid );
  input [31:0] N_RxData;
  input [31:0] S_RxData;
  input [31:0] W_RxData;
  input [31:0] E_RxData;
  input [31:0] Packet_From_Node;
  output [31:0] N_TxData;
  output [31:0] S_TxData;
  output [31:0] W_TxData;
  output [31:0] E_TxData;
  output [31:0] Packet_To_Node;
  input Clk_r, Rst_n, N_Tx_Ready, N_Tx_Error, N_RxData_Valid, S_Tx_Ready,
         S_Tx_Error, S_RxData_Valid, W_Tx_Ready, W_Tx_Error, W_RxData_Valid,
         E_Tx_Ready, E_Tx_Error, E_RxData_Valid, Packet_From_Node_Valid;
  output N_TxData_Valid, N_Error_Ack, N_Core_Rcv_Ready, S_TxData_Valid,
         S_Error_Ack, S_Core_Rcv_Ready, W_TxData_Valid, W_Error_Ack,
         W_Core_Rcv_Ready, E_TxData_Valid, E_Error_Ack, E_Core_Rcv_Ready,
         Core_Load_Ack, Packet_To_Node_Valid;
  wire   N_TxQueue_Write, N_RxQueue_Read, N_RxQueue_Empty, N_TxQueue_Full,
         S_TxQueue_Write, S_RxQueue_Read, S_RxQueue_Empty, S_TxQueue_Full,
         E_TxQueue_Write, E_RxQueue_Read, E_RxQueue_Empty, E_TxQueue_Full,
         W_TxQueue_Write, W_RxQueue_Read, W_RxQueue_Empty, W_TxQueue_Full,
         NM_Empty, NM_Full, NM_Read, NM_Write;
  wire   [31:0] N_Tx_Packet;
  wire   [31:0] N_Rx_Packet;
  wire   [31:0] S_Tx_Packet;
  wire   [31:0] S_Rx_Packet;
  wire   [31:0] E_Tx_Packet;
  wire   [31:0] E_Rx_Packet;
  wire   [31:0] W_Tx_Packet;
  wire   [31:0] W_Rx_Packet;
  wire   [7:0] Router_Addr;
  wire   [3:0] Link_Config;
  wire   [31:0] NM_In_Packet;
  wire   [31:0] NM_Out_Packet;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7;

  Link_Control_0 N_Link_Control ( .Clk_r(Clk_r), .Rst_n(Rst_n), .Tx_Ready(
        N_Tx_Ready), .Tx_Error(N_Tx_Error), .RxData_Valid(N_RxData_Valid), 
        .RxData(N_RxData), .Packet_From_Core(N_Tx_Packet), .TxQueue_Write(
        N_TxQueue_Write), .RxQueue_Read(N_RxQueue_Read), .TxData_Valid(
        N_TxData_Valid), .TxData(N_TxData), .Error_Ack(N_Error_Ack), 
        .Core_Rcv_Ready(N_Core_Rcv_Ready), .Packet_To_Core(N_Rx_Packet), 
        .RxQueue_Empty(N_RxQueue_Empty), .TxQueue_Full(N_TxQueue_Full) );
  Link_Control_3 S_Link_Control ( .Clk_r(Clk_r), .Rst_n(Rst_n), .Tx_Ready(
        S_Tx_Ready), .Tx_Error(S_Tx_Error), .RxData_Valid(S_RxData_Valid), 
        .RxData(S_RxData), .Packet_From_Core(S_Tx_Packet), .TxQueue_Write(
        S_TxQueue_Write), .RxQueue_Read(S_RxQueue_Read), .TxData_Valid(
        S_TxData_Valid), .TxData(S_TxData), .Error_Ack(S_Error_Ack), 
        .Core_Rcv_Ready(S_Core_Rcv_Ready), .Packet_To_Core(S_Rx_Packet), 
        .RxQueue_Empty(S_RxQueue_Empty), .TxQueue_Full(S_TxQueue_Full) );
  Link_Control_2 E_Link_Control ( .Clk_r(Clk_r), .Rst_n(Rst_n), .Tx_Ready(
        E_Tx_Ready), .Tx_Error(E_Tx_Error), .RxData_Valid(E_RxData_Valid), 
        .RxData(E_RxData), .Packet_From_Core(E_Tx_Packet), .TxQueue_Write(
        E_TxQueue_Write), .RxQueue_Read(E_RxQueue_Read), .TxData_Valid(
        E_TxData_Valid), .TxData(E_TxData), .Error_Ack(E_Error_Ack), 
        .Core_Rcv_Ready(E_Core_Rcv_Ready), .Packet_To_Core(E_Rx_Packet), 
        .RxQueue_Empty(E_RxQueue_Empty), .TxQueue_Full(E_TxQueue_Full) );
  Link_Control_1 W_Link_Control ( .Clk_r(Clk_r), .Rst_n(Rst_n), .Tx_Ready(
        W_Tx_Ready), .Tx_Error(W_Tx_Error), .RxData_Valid(W_RxData_Valid), 
        .RxData(W_RxData), .Packet_From_Core(W_Tx_Packet), .TxQueue_Write(
        W_TxQueue_Write), .RxQueue_Read(W_RxQueue_Read), .TxData_Valid(
        W_TxData_Valid), .TxData(W_TxData), .Error_Ack(W_Error_Ack), 
        .Core_Rcv_Ready(W_Core_Rcv_Ready), .Packet_To_Core(W_Rx_Packet), 
        .RxQueue_Empty(W_RxQueue_Empty), .TxQueue_Full(W_TxQueue_Full) );
  Routing_State_Machine routing_state_machine ( .Clk_r(Clk_r), .Rst_n(Rst_n), 
        .Router_Address(Router_Addr), .Link_Config(Link_Config), 
        .Packet_From_Link_N(N_Rx_Packet), .Packet_From_Link_S(S_Rx_Packet), 
        .Packet_From_Link_W(W_Rx_Packet), .Packet_From_Link_E(E_Rx_Packet), 
        .Packet_From_Node({NM_In_Packet[31:24], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, NM_In_Packet[15:0]}), .RxQueue_Empty_N(
        N_RxQueue_Empty), .RxQueue_Empty_S(S_RxQueue_Empty), .RxQueue_Empty_W(
        W_RxQueue_Empty), .RxQueue_Empty_E(E_RxQueue_Empty), .TxQueue_Full_N(
        N_TxQueue_Full), .TxQueue_Full_S(S_TxQueue_Full), .TxQueue_Full_W(
        W_TxQueue_Full), .TxQueue_Full_E(E_TxQueue_Full), .To_Node_Full(
        NM_Full), .Node_Queue_Empty(NM_Empty), .Packet_To_Link_N(N_Tx_Packet), 
        .Packet_To_Link_S(S_Tx_Packet), .Packet_To_Link_W(W_Tx_Packet), 
        .Packet_To_Link_E(E_Tx_Packet), .Packet_To_Node(NM_Out_Packet), 
        .TxQueue_Write_N(N_TxQueue_Write), .TxQueue_Write_S(S_TxQueue_Write), 
        .TxQueue_Write_W(W_TxQueue_Write), .TxQueue_Write_E(E_TxQueue_Write), 
        .To_Node_Write(NM_Write), .RxQueue_Read_N(N_RxQueue_Read), 
        .RxQueue_Read_S(S_RxQueue_Read), .RxQueue_Read_W(W_RxQueue_Read), 
        .RxQueue_Read_E(E_RxQueue_Read), .Node_Read(NM_Read) );
  Node_Manager node_manager ( .Clk_r(Clk_r), .Rst_n(Rst_n), .Packet_From_Core(
        NM_Out_Packet), .Packet_From_Node(Packet_From_Node), 
        .Packet_From_Node_Valid(Packet_From_Node_Valid), .Read_Packet(NM_Read), 
        .To_Node_Write(NM_Write), .Router_Address(Router_Addr), .Link_Config(
        Link_Config), .Packet_To_Core({NM_In_Packet[31:24], 
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, NM_In_Packet[15:0]}), 
        .Packet_To_Node(Packet_To_Node), .Packet_To_Node_Valid(
        Packet_To_Node_Valid), .Core_Load_Ack(Core_Load_Ack), .Queue_Empty(
        NM_Empty), .To_Node_Full(NM_Full) );
endmodule

