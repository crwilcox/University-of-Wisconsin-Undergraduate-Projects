library verilog;
use verilog.vl_types.all;
entity p1_mealy_tb is
end p1_mealy_tb;
