library verilog;
use verilog.vl_types.all;
entity register_file_16_tb is
end register_file_16_tb;
