library verilog;
use verilog.vl_types.all;
entity decoder_2_to_4_139 is
    port(
        E               : in     vl_logic;
        A0              : in     vl_logic;
        A1              : in     vl_logic;
        O0              : out    vl_logic;
        O1              : out    vl_logic;
        O2              : out    vl_logic;
        O3              : out    vl_logic
    );
end decoder_2_to_4_139;
