library verilog;
use verilog.vl_types.all;
entity p2_tb is
end p2_tb;
