
module Packet_Queue_synth ( Clk_r, Rst_n, Packet_In, Read_Ack, Write_Ack, Packet_Out, 
        Empty, Full );
  input [31:0] Packet_In;
  output [31:0] Packet_Out;
  input Clk_r, Rst_n, Read_Ack, Write_Ack;
  output Empty, Full;
  wire   \Queue[4][31] , \Queue[4][30] , \Queue[4][29] , \Queue[4][28] ,
         \Queue[4][27] , \Queue[4][26] , \Queue[4][25] , \Queue[4][24] ,
         \Queue[4][23] , \Queue[4][22] , \Queue[4][21] , \Queue[4][20] ,
         \Queue[4][19] , \Queue[4][18] , \Queue[4][17] , \Queue[4][16] ,
         \Queue[4][15] , \Queue[4][14] , \Queue[4][13] , \Queue[4][12] ,
         \Queue[4][11] , \Queue[4][10] , \Queue[4][9] , \Queue[4][8] ,
         \Queue[4][7] , \Queue[4][6] , \Queue[4][5] , \Queue[4][4] ,
         \Queue[4][3] , \Queue[4][2] , \Queue[4][1] , \Queue[4][0] ,
         \Queue[3][31] , \Queue[3][30] , \Queue[3][29] , \Queue[3][28] ,
         \Queue[3][27] , \Queue[3][26] , \Queue[3][25] , \Queue[3][24] ,
         \Queue[3][23] , \Queue[3][22] , \Queue[3][21] , \Queue[3][20] ,
         \Queue[3][19] , \Queue[3][18] , \Queue[3][17] , \Queue[3][16] ,
         \Queue[3][15] , \Queue[3][14] , \Queue[3][13] , \Queue[3][12] ,
         \Queue[3][11] , \Queue[3][10] , \Queue[3][9] , \Queue[3][8] ,
         \Queue[3][7] , \Queue[3][6] , \Queue[3][5] , \Queue[3][4] ,
         \Queue[3][3] , \Queue[3][2] , \Queue[3][1] , \Queue[3][0] ,
         \Queue[2][31] , \Queue[2][30] , \Queue[2][29] , \Queue[2][28] ,
         \Queue[2][27] , \Queue[2][26] , \Queue[2][25] , \Queue[2][24] ,
         \Queue[2][23] , \Queue[2][22] , \Queue[2][21] , \Queue[2][20] ,
         \Queue[2][19] , \Queue[2][18] , \Queue[2][17] , \Queue[2][16] ,
         \Queue[2][15] , \Queue[2][14] , \Queue[2][13] , \Queue[2][12] ,
         \Queue[2][11] , \Queue[2][10] , \Queue[2][9] , \Queue[2][8] ,
         \Queue[2][7] , \Queue[2][6] , \Queue[2][5] , \Queue[2][4] ,
         \Queue[2][3] , \Queue[2][2] , \Queue[2][1] , \Queue[2][0] ,
         \Queue[1][31] , \Queue[1][30] , \Queue[1][29] , \Queue[1][28] ,
         \Queue[1][27] , \Queue[1][26] , \Queue[1][25] , \Queue[1][24] ,
         \Queue[1][23] , \Queue[1][22] , \Queue[1][21] , \Queue[1][20] ,
         \Queue[1][19] , \Queue[1][18] , \Queue[1][17] , \Queue[1][16] ,
         \Queue[1][15] , \Queue[1][14] , \Queue[1][13] , \Queue[1][12] ,
         \Queue[1][11] , \Queue[1][10] , \Queue[1][9] , \Queue[1][8] ,
         \Queue[1][7] , \Queue[1][6] , \Queue[1][5] , \Queue[1][4] ,
         \Queue[1][3] , \Queue[1][2] , \Queue[1][1] , \Queue[1][0] , n1, n2,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574;
  wire   [2:0] Count;

  FDN1QM1P \Queue_reg[4][30]  ( .D(n338), .CPN(Clk_r), .Q(\Queue[4][30] ) );
  FDN1QM1P \Queue_reg[3][30]  ( .D(n210), .CPN(Clk_r), .Q(\Queue[3][30] ) );
  FDN1QM1P \Queue_reg[2][30]  ( .D(n242), .CPN(Clk_r), .Q(\Queue[2][30] ) );
  FDN1QM1P \Queue_reg[4][29]  ( .D(n339), .CPN(Clk_r), .Q(\Queue[4][29] ) );
  FDN1QM1P \Queue_reg[3][29]  ( .D(n211), .CPN(Clk_r), .Q(\Queue[3][29] ) );
  FDN1QM1P \Queue_reg[2][29]  ( .D(n243), .CPN(Clk_r), .Q(\Queue[2][29] ) );
  FDN1QM1P \Queue_reg[4][28]  ( .D(n340), .CPN(Clk_r), .Q(\Queue[4][28] ) );
  FDN1QM1P \Queue_reg[3][28]  ( .D(n212), .CPN(Clk_r), .Q(\Queue[3][28] ) );
  FDN1QM1P \Queue_reg[2][28]  ( .D(n244), .CPN(Clk_r), .Q(\Queue[2][28] ) );
  FDN1QM1P \Queue_reg[4][27]  ( .D(n341), .CPN(Clk_r), .Q(\Queue[4][27] ) );
  FDN1QM1P \Queue_reg[3][27]  ( .D(n213), .CPN(Clk_r), .Q(\Queue[3][27] ) );
  FDN1QM1P \Queue_reg[2][27]  ( .D(n245), .CPN(Clk_r), .Q(\Queue[2][27] ) );
  FDN1QM1P \Queue_reg[4][26]  ( .D(n342), .CPN(Clk_r), .Q(\Queue[4][26] ) );
  FDN1QM1P \Queue_reg[3][26]  ( .D(n214), .CPN(Clk_r), .Q(\Queue[3][26] ) );
  FDN1QM1P \Queue_reg[2][26]  ( .D(n246), .CPN(Clk_r), .Q(\Queue[2][26] ) );
  FDN1QM1P \Queue_reg[4][25]  ( .D(n343), .CPN(Clk_r), .Q(\Queue[4][25] ) );
  FDN1QM1P \Queue_reg[3][25]  ( .D(n215), .CPN(Clk_r), .Q(\Queue[3][25] ) );
  FDN1QM1P \Queue_reg[2][25]  ( .D(n247), .CPN(Clk_r), .Q(\Queue[2][25] ) );
  FDN1QM1P \Queue_reg[4][24]  ( .D(n344), .CPN(Clk_r), .Q(\Queue[4][24] ) );
  FDN1QM1P \Queue_reg[3][24]  ( .D(n216), .CPN(Clk_r), .Q(\Queue[3][24] ) );
  FDN1QM1P \Queue_reg[2][24]  ( .D(n248), .CPN(Clk_r), .Q(\Queue[2][24] ) );
  FDN1QM1P \Queue_reg[4][23]  ( .D(n345), .CPN(Clk_r), .Q(\Queue[4][23] ) );
  FDN1QM1P \Queue_reg[3][23]  ( .D(n217), .CPN(Clk_r), .Q(\Queue[3][23] ) );
  FDN1QM1P \Queue_reg[2][23]  ( .D(n249), .CPN(Clk_r), .Q(\Queue[2][23] ) );
  FDN1QM1P \Queue_reg[4][22]  ( .D(n346), .CPN(Clk_r), .Q(\Queue[4][22] ) );
  FDN1QM1P \Queue_reg[3][22]  ( .D(n218), .CPN(Clk_r), .Q(\Queue[3][22] ) );
  FDN1QM1P \Queue_reg[2][22]  ( .D(n250), .CPN(Clk_r), .Q(\Queue[2][22] ) );
  FDN1QM1P \Queue_reg[4][21]  ( .D(n347), .CPN(Clk_r), .Q(\Queue[4][21] ) );
  FDN1QM1P \Queue_reg[3][21]  ( .D(n219), .CPN(Clk_r), .Q(\Queue[3][21] ) );
  FDN1QM1P \Queue_reg[2][21]  ( .D(n251), .CPN(Clk_r), .Q(\Queue[2][21] ) );
  FDN1QM1P \Queue_reg[4][20]  ( .D(n348), .CPN(Clk_r), .Q(\Queue[4][20] ) );
  FDN1QM1P \Queue_reg[3][20]  ( .D(n220), .CPN(Clk_r), .Q(\Queue[3][20] ) );
  FDN1QM1P \Queue_reg[2][20]  ( .D(n252), .CPN(Clk_r), .Q(\Queue[2][20] ) );
  FDN1QM1P \Queue_reg[4][19]  ( .D(n349), .CPN(Clk_r), .Q(\Queue[4][19] ) );
  FDN1QM1P \Queue_reg[3][19]  ( .D(n221), .CPN(Clk_r), .Q(\Queue[3][19] ) );
  FDN1QM1P \Queue_reg[2][19]  ( .D(n253), .CPN(Clk_r), .Q(\Queue[2][19] ) );
  FDN1QM1P \Queue_reg[4][18]  ( .D(n350), .CPN(Clk_r), .Q(\Queue[4][18] ) );
  FDN1QM1P \Queue_reg[3][18]  ( .D(n222), .CPN(Clk_r), .Q(\Queue[3][18] ) );
  FDN1QM1P \Queue_reg[2][18]  ( .D(n254), .CPN(Clk_r), .Q(\Queue[2][18] ) );
  FDN1QM1P \Queue_reg[4][17]  ( .D(n351), .CPN(Clk_r), .Q(\Queue[4][17] ) );
  FDN1QM1P \Queue_reg[3][17]  ( .D(n223), .CPN(Clk_r), .Q(\Queue[3][17] ) );
  FDN1QM1P \Queue_reg[2][17]  ( .D(n255), .CPN(Clk_r), .Q(\Queue[2][17] ) );
  FDN1QM1P \Queue_reg[4][16]  ( .D(n352), .CPN(Clk_r), .Q(\Queue[4][16] ) );
  FDN1QM1P \Queue_reg[3][16]  ( .D(n224), .CPN(Clk_r), .Q(\Queue[3][16] ) );
  FDN1QM1P \Queue_reg[2][16]  ( .D(n256), .CPN(Clk_r), .Q(\Queue[2][16] ) );
  FDN1QM1P \Queue_reg[4][15]  ( .D(n353), .CPN(Clk_r), .Q(\Queue[4][15] ) );
  FDN1QM1P \Queue_reg[3][15]  ( .D(n225), .CPN(Clk_r), .Q(\Queue[3][15] ) );
  FDN1QM1P \Queue_reg[2][15]  ( .D(n257), .CPN(Clk_r), .Q(\Queue[2][15] ) );
  FDN1QM1P \Queue_reg[4][14]  ( .D(n354), .CPN(Clk_r), .Q(\Queue[4][14] ) );
  FDN1QM1P \Queue_reg[3][14]  ( .D(n226), .CPN(Clk_r), .Q(\Queue[3][14] ) );
  FDN1QM1P \Queue_reg[2][14]  ( .D(n258), .CPN(Clk_r), .Q(\Queue[2][14] ) );
  FDN1QM1P \Queue_reg[4][13]  ( .D(n355), .CPN(Clk_r), .Q(\Queue[4][13] ) );
  FDN1QM1P \Queue_reg[3][13]  ( .D(n227), .CPN(Clk_r), .Q(\Queue[3][13] ) );
  FDN1QM1P \Queue_reg[2][13]  ( .D(n259), .CPN(Clk_r), .Q(\Queue[2][13] ) );
  FDN1QM1P \Queue_reg[4][12]  ( .D(n356), .CPN(Clk_r), .Q(\Queue[4][12] ) );
  FDN1QM1P \Queue_reg[3][12]  ( .D(n228), .CPN(Clk_r), .Q(\Queue[3][12] ) );
  FDN1QM1P \Queue_reg[2][12]  ( .D(n260), .CPN(Clk_r), .Q(\Queue[2][12] ) );
  FDN1QM1P \Queue_reg[4][11]  ( .D(n357), .CPN(Clk_r), .Q(\Queue[4][11] ) );
  FDN1QM1P \Queue_reg[3][11]  ( .D(n229), .CPN(Clk_r), .Q(\Queue[3][11] ) );
  FDN1QM1P \Queue_reg[2][11]  ( .D(n261), .CPN(Clk_r), .Q(\Queue[2][11] ) );
  FDN1QM1P \Queue_reg[4][10]  ( .D(n358), .CPN(Clk_r), .Q(\Queue[4][10] ) );
  FDN1QM1P \Queue_reg[3][10]  ( .D(n230), .CPN(Clk_r), .Q(\Queue[3][10] ) );
  FDN1QM1P \Queue_reg[2][10]  ( .D(n262), .CPN(Clk_r), .Q(\Queue[2][10] ) );
  FDN1QM1P \Queue_reg[4][9]  ( .D(n359), .CPN(Clk_r), .Q(\Queue[4][9] ) );
  FDN1QM1P \Queue_reg[3][9]  ( .D(n231), .CPN(Clk_r), .Q(\Queue[3][9] ) );
  FDN1QM1P \Queue_reg[2][9]  ( .D(n263), .CPN(Clk_r), .Q(\Queue[2][9] ) );
  FDN1QM1P \Queue_reg[4][8]  ( .D(n360), .CPN(Clk_r), .Q(\Queue[4][8] ) );
  FDN1QM1P \Queue_reg[3][8]  ( .D(n232), .CPN(Clk_r), .Q(\Queue[3][8] ) );
  FDN1QM1P \Queue_reg[2][8]  ( .D(n264), .CPN(Clk_r), .Q(\Queue[2][8] ) );
  FDN1QM1P \Queue_reg[4][7]  ( .D(n361), .CPN(Clk_r), .Q(\Queue[4][7] ) );
  FDN1QM1P \Queue_reg[3][7]  ( .D(n233), .CPN(Clk_r), .Q(\Queue[3][7] ) );
  FDN1QM1P \Queue_reg[2][7]  ( .D(n265), .CPN(Clk_r), .Q(\Queue[2][7] ) );
  FDN1QM1P \Queue_reg[4][6]  ( .D(n362), .CPN(Clk_r), .Q(\Queue[4][6] ) );
  FDN1QM1P \Queue_reg[3][6]  ( .D(n234), .CPN(Clk_r), .Q(\Queue[3][6] ) );
  FDN1QM1P \Queue_reg[2][6]  ( .D(n266), .CPN(Clk_r), .Q(\Queue[2][6] ) );
  FDN1QM1P \Queue_reg[4][5]  ( .D(n363), .CPN(Clk_r), .Q(\Queue[4][5] ) );
  FDN1QM1P \Queue_reg[3][5]  ( .D(n235), .CPN(Clk_r), .Q(\Queue[3][5] ) );
  FDN1QM1P \Queue_reg[2][5]  ( .D(n267), .CPN(Clk_r), .Q(\Queue[2][5] ) );
  FDN1QM1P \Queue_reg[4][4]  ( .D(n364), .CPN(Clk_r), .Q(\Queue[4][4] ) );
  FDN1QM1P \Queue_reg[3][4]  ( .D(n236), .CPN(Clk_r), .Q(\Queue[3][4] ) );
  FDN1QM1P \Queue_reg[2][4]  ( .D(n268), .CPN(Clk_r), .Q(\Queue[2][4] ) );
  FDN1QM1P \Queue_reg[4][3]  ( .D(n365), .CPN(Clk_r), .Q(\Queue[4][3] ) );
  FDN1QM1P \Queue_reg[3][3]  ( .D(n237), .CPN(Clk_r), .Q(\Queue[3][3] ) );
  FDN1QM1P \Queue_reg[2][3]  ( .D(n269), .CPN(Clk_r), .Q(\Queue[2][3] ) );
  FDN1QM1P \Queue_reg[4][2]  ( .D(n366), .CPN(Clk_r), .Q(\Queue[4][2] ) );
  FDN1QM1P \Queue_reg[3][2]  ( .D(n238), .CPN(Clk_r), .Q(\Queue[3][2] ) );
  FDN1QM1P \Queue_reg[2][2]  ( .D(n270), .CPN(Clk_r), .Q(\Queue[2][2] ) );
  FDN1QM1P \Queue_reg[4][1]  ( .D(n367), .CPN(Clk_r), .Q(\Queue[4][1] ) );
  FDN1QM1P \Queue_reg[3][1]  ( .D(n239), .CPN(Clk_r), .Q(\Queue[3][1] ) );
  FDN1QM1P \Queue_reg[2][1]  ( .D(n271), .CPN(Clk_r), .Q(\Queue[2][1] ) );
  FDN1QM1P \Queue_reg[4][0]  ( .D(n368), .CPN(Clk_r), .Q(\Queue[4][0] ) );
  FDN1QM1P \Queue_reg[3][0]  ( .D(n240), .CPN(Clk_r), .Q(\Queue[3][0] ) );
  FDN1QM1P \Queue_reg[2][0]  ( .D(n272), .CPN(Clk_r), .Q(\Queue[2][0] ) );
  FDN1QM1P \Queue_reg[4][31]  ( .D(n369), .CPN(Clk_r), .Q(\Queue[4][31] ) );
  FDN1QM1P \Queue_reg[3][31]  ( .D(n209), .CPN(Clk_r), .Q(\Queue[3][31] ) );
  FDN1QM1P \Queue_reg[2][31]  ( .D(n241), .CPN(Clk_r), .Q(\Queue[2][31] ) );
  FDN1QM1P \Queue_reg[1][31]  ( .D(n305), .CPN(Clk_r), .Q(\Queue[1][31] ) );
  FDN1QM1P \Queue_reg[0][31]  ( .D(n273), .CPN(Clk_r), .Q(Packet_Out[31]) );
  FDN1QM1P \Queue_reg[1][30]  ( .D(n306), .CPN(Clk_r), .Q(\Queue[1][30] ) );
  FDN1QM1P \Queue_reg[0][30]  ( .D(n274), .CPN(Clk_r), .Q(Packet_Out[30]) );
  FDN1QM1P \Queue_reg[1][29]  ( .D(n307), .CPN(Clk_r), .Q(\Queue[1][29] ) );
  FDN1QM1P \Queue_reg[0][29]  ( .D(n275), .CPN(Clk_r), .Q(Packet_Out[29]) );
  FDN1QM1P \Queue_reg[1][28]  ( .D(n308), .CPN(Clk_r), .Q(\Queue[1][28] ) );
  FDN1QM1P \Queue_reg[0][28]  ( .D(n276), .CPN(Clk_r), .Q(Packet_Out[28]) );
  FDN1QM1P \Queue_reg[1][27]  ( .D(n309), .CPN(Clk_r), .Q(\Queue[1][27] ) );
  FDN1QM1P \Queue_reg[0][27]  ( .D(n277), .CPN(Clk_r), .Q(Packet_Out[27]) );
  FDN1QM1P \Queue_reg[1][26]  ( .D(n310), .CPN(Clk_r), .Q(\Queue[1][26] ) );
  FDN1QM1P \Queue_reg[0][26]  ( .D(n278), .CPN(Clk_r), .Q(Packet_Out[26]) );
  FDN1QM1P \Queue_reg[1][25]  ( .D(n311), .CPN(Clk_r), .Q(\Queue[1][25] ) );
  FDN1QM1P \Queue_reg[0][25]  ( .D(n279), .CPN(Clk_r), .Q(Packet_Out[25]) );
  FDN1QM1P \Queue_reg[1][24]  ( .D(n312), .CPN(Clk_r), .Q(\Queue[1][24] ) );
  FDN1QM1P \Queue_reg[0][24]  ( .D(n280), .CPN(Clk_r), .Q(Packet_Out[24]) );
  FDN1QM1P \Queue_reg[1][23]  ( .D(n313), .CPN(Clk_r), .Q(\Queue[1][23] ) );
  FDN1QM1P \Queue_reg[0][23]  ( .D(n281), .CPN(Clk_r), .Q(Packet_Out[23]) );
  FDN1QM1P \Queue_reg[1][22]  ( .D(n314), .CPN(Clk_r), .Q(\Queue[1][22] ) );
  FDN1QM1P \Queue_reg[0][22]  ( .D(n282), .CPN(Clk_r), .Q(Packet_Out[22]) );
  FDN1QM1P \Queue_reg[1][21]  ( .D(n315), .CPN(Clk_r), .Q(\Queue[1][21] ) );
  FDN1QM1P \Queue_reg[0][21]  ( .D(n283), .CPN(Clk_r), .Q(Packet_Out[21]) );
  FDN1QM1P \Queue_reg[1][20]  ( .D(n316), .CPN(Clk_r), .Q(\Queue[1][20] ) );
  FDN1QM1P \Queue_reg[0][20]  ( .D(n284), .CPN(Clk_r), .Q(Packet_Out[20]) );
  FDN1QM1P \Queue_reg[1][19]  ( .D(n317), .CPN(Clk_r), .Q(\Queue[1][19] ) );
  FDN1QM1P \Queue_reg[0][19]  ( .D(n285), .CPN(Clk_r), .Q(Packet_Out[19]) );
  FDN1QM1P \Queue_reg[1][18]  ( .D(n318), .CPN(Clk_r), .Q(\Queue[1][18] ) );
  FDN1QM1P \Queue_reg[0][18]  ( .D(n286), .CPN(Clk_r), .Q(Packet_Out[18]) );
  FDN1QM1P \Queue_reg[1][17]  ( .D(n319), .CPN(Clk_r), .Q(\Queue[1][17] ) );
  FDN1QM1P \Queue_reg[0][17]  ( .D(n287), .CPN(Clk_r), .Q(Packet_Out[17]) );
  FDN1QM1P \Queue_reg[1][16]  ( .D(n320), .CPN(Clk_r), .Q(\Queue[1][16] ) );
  FDN1QM1P \Queue_reg[0][16]  ( .D(n288), .CPN(Clk_r), .Q(Packet_Out[16]) );
  FDN1QM1P \Queue_reg[1][15]  ( .D(n321), .CPN(Clk_r), .Q(\Queue[1][15] ) );
  FDN1QM1P \Queue_reg[0][15]  ( .D(n289), .CPN(Clk_r), .Q(Packet_Out[15]) );
  FDN1QM1P \Queue_reg[1][14]  ( .D(n322), .CPN(Clk_r), .Q(\Queue[1][14] ) );
  FDN1QM1P \Queue_reg[0][14]  ( .D(n290), .CPN(Clk_r), .Q(Packet_Out[14]) );
  FDN1QM1P \Queue_reg[1][13]  ( .D(n323), .CPN(Clk_r), .Q(\Queue[1][13] ) );
  FDN1QM1P \Queue_reg[0][13]  ( .D(n291), .CPN(Clk_r), .Q(Packet_Out[13]) );
  FDN1QM1P \Queue_reg[1][12]  ( .D(n324), .CPN(Clk_r), .Q(\Queue[1][12] ) );
  FDN1QM1P \Queue_reg[0][12]  ( .D(n292), .CPN(Clk_r), .Q(Packet_Out[12]) );
  FDN1QM1P \Queue_reg[1][11]  ( .D(n325), .CPN(Clk_r), .Q(\Queue[1][11] ) );
  FDN1QM1P \Queue_reg[0][11]  ( .D(n293), .CPN(Clk_r), .Q(Packet_Out[11]) );
  FDN1QM1P \Queue_reg[1][10]  ( .D(n326), .CPN(Clk_r), .Q(\Queue[1][10] ) );
  FDN1QM1P \Queue_reg[0][10]  ( .D(n294), .CPN(Clk_r), .Q(Packet_Out[10]) );
  FDN1QM1P \Queue_reg[1][9]  ( .D(n327), .CPN(Clk_r), .Q(\Queue[1][9] ) );
  FDN1QM1P \Queue_reg[0][9]  ( .D(n295), .CPN(Clk_r), .Q(Packet_Out[9]) );
  FDN1QM1P \Queue_reg[1][8]  ( .D(n328), .CPN(Clk_r), .Q(\Queue[1][8] ) );
  FDN1QM1P \Queue_reg[0][8]  ( .D(n296), .CPN(Clk_r), .Q(Packet_Out[8]) );
  FDN1QM1P \Queue_reg[1][7]  ( .D(n329), .CPN(Clk_r), .Q(\Queue[1][7] ) );
  FDN1QM1P \Queue_reg[0][7]  ( .D(n297), .CPN(Clk_r), .Q(Packet_Out[7]) );
  FDN1QM1P \Queue_reg[1][6]  ( .D(n330), .CPN(Clk_r), .Q(\Queue[1][6] ) );
  FDN1QM1P \Queue_reg[0][6]  ( .D(n298), .CPN(Clk_r), .Q(Packet_Out[6]) );
  FDN1QM1P \Queue_reg[1][5]  ( .D(n331), .CPN(Clk_r), .Q(\Queue[1][5] ) );
  FDN1QM1P \Queue_reg[0][5]  ( .D(n299), .CPN(Clk_r), .Q(Packet_Out[5]) );
  FDN1QM1P \Queue_reg[1][4]  ( .D(n332), .CPN(Clk_r), .Q(\Queue[1][4] ) );
  FDN1QM1P \Queue_reg[0][4]  ( .D(n300), .CPN(Clk_r), .Q(Packet_Out[4]) );
  FDN1QM1P \Queue_reg[1][3]  ( .D(n333), .CPN(Clk_r), .Q(\Queue[1][3] ) );
  FDN1QM1P \Queue_reg[0][3]  ( .D(n301), .CPN(Clk_r), .Q(Packet_Out[3]) );
  FDN1QM1P \Queue_reg[1][2]  ( .D(n334), .CPN(Clk_r), .Q(\Queue[1][2] ) );
  FDN1QM1P \Queue_reg[0][2]  ( .D(n302), .CPN(Clk_r), .Q(Packet_Out[2]) );
  FDN1QM1P \Queue_reg[1][1]  ( .D(n335), .CPN(Clk_r), .Q(\Queue[1][1] ) );
  FDN1QM1P \Queue_reg[0][1]  ( .D(n303), .CPN(Clk_r), .Q(Packet_Out[1]) );
  FDN1QM1P \Queue_reg[1][0]  ( .D(n336), .CPN(Clk_r), .Q(\Queue[1][0] ) );
  FDN1QM1P \Queue_reg[0][0]  ( .D(n304), .CPN(Clk_r), .Q(Packet_Out[0]) );
  FDN2QM1P Empty_reg ( .D(n1), .CPN(Clk_r), .CD(Rst_n), .Q(n2) );
  FDN2QM1P Full_reg ( .D(n337), .CPN(Clk_r), .CD(Rst_n), .Q(Full) );
  FDN2QM1P \Count_reg[0]  ( .D(n372), .CPN(Clk_r), .CD(Rst_n), .Q(Count[0]) );
  FDN2QM1P \Count_reg[1]  ( .D(n371), .CPN(Clk_r), .CD(Rst_n), .Q(Count[1]) );
  FDN2QM1P \Count_reg[2]  ( .D(n370), .CPN(Clk_r), .CD(Rst_n), .Q(Count[2]) );
  N1M1P U375 ( .A(Count[2]), .Z(n393) );
  NR3M1P U376 ( .A(Count[0]), .B(Count[1]), .C(n393), .Z(n507) );
  OAI211M4P U377 ( .A(n574), .B(n502), .C(Write_Ack), .D(n432), .Z(n376) );
  N1M3P U378 ( .A(n384), .Z(n385) );
  OAI211M4P U379 ( .A(n468), .B(n504), .C(Rst_n), .D(n503), .Z(n375) );
  OAI211M4P U380 ( .A(n505), .B(n504), .C(Rst_n), .D(n503), .Z(n382) );
  OAI211M4P U381 ( .A(n507), .B(n502), .C(Write_Ack), .D(n501), .Z(n377) );
  NR2I1M8P U382 ( .A(n431), .B(n394), .Z(n383) );
  OAI211M4P U383 ( .A(n505), .B(n502), .C(Write_Ack), .D(n466), .Z(n373) );
  OAI211M4P U384 ( .A(n468), .B(n502), .C(Write_Ack), .D(n397), .Z(n374) );
  N1M1P U385 ( .A(n432), .Z(n464) );
  AND3M1P U386 ( .A(n393), .B(Count[0]), .C(Count[1]), .Z(n505) );
  N1M1P U387 ( .A(Count[1]), .Z(n395) );
  N1M1P U388 ( .A(Count[0]), .Z(n396) );
  N1M1P U389 ( .A(Write_Ack), .Z(n467) );
  OA21M1P U390 ( .A(Write_Ack), .B(Read_Ack), .C(n397), .Z(n384) );
  AOI21M6P U391 ( .A(Write_Ack), .B(n468), .C(n506), .Z(n378) );
  N1M1P U392 ( .A(n507), .Z(n394) );
  AOI21M6P U393 ( .A(Write_Ack), .B(n505), .C(n506), .Z(n380) );
  AOI21M6P U394 ( .A(Write_Ack), .B(n574), .C(n506), .Z(n379) );
  AOI21M6P U395 ( .A(Write_Ack), .B(n507), .C(n506), .Z(n381) );
  AND3M1P U396 ( .A(Count[0]), .B(n393), .C(n395), .Z(n574) );
  N1M2P U397 ( .A(n392), .Z(n504) );
  N1M2P U398 ( .A(n432), .Z(n386) );
  NR2M2P U399 ( .A(Read_Ack), .B(n467), .Z(n392) );
  NR3M2P U400 ( .A(Count[0]), .B(Count[2]), .C(n395), .Z(n468) );
  OAI21M1P U401 ( .A(n431), .B(n430), .C(n506), .Z(n432) );
  ND3M1P U402 ( .A(n396), .B(n393), .C(n395), .Z(n430) );
  N1M1P U403 ( .A(Read_Ack), .Z(n502) );
  ND2M1P U404 ( .A(Read_Ack), .B(Rst_n), .Z(n506) );
  ND2M1P U405 ( .A(n392), .B(Rst_n), .Z(n431) );
  N1M1P U406 ( .A(Packet_In[8]), .Z(n525) );
  N1M1P U407 ( .A(Packet_In[12]), .Z(n533) );
  N1M1P U408 ( .A(Packet_In[25]), .Z(n559) );
  N1M1P U409 ( .A(Packet_In[24]), .Z(n557) );
  N1M1P U410 ( .A(Packet_In[14]), .Z(n537) );
  N1M1P U411 ( .A(Packet_In[17]), .Z(n543) );
  N1M1P U412 ( .A(Packet_In[16]), .Z(n541) );
  N1M1P U413 ( .A(Packet_In[30]), .Z(n569) );
  N1M1P U414 ( .A(Packet_In[27]), .Z(n563) );
  N1M1P U415 ( .A(Packet_In[31]), .Z(n571) );
  N1M1P U416 ( .A(Packet_In[0]), .Z(n509) );
  N1M1P U417 ( .A(Packet_In[5]), .Z(n519) );
  N1M1P U418 ( .A(Packet_In[2]), .Z(n513) );
  N1M1P U419 ( .A(Packet_In[15]), .Z(n539) );
  N1M1P U420 ( .A(Packet_In[3]), .Z(n515) );
  N1M1P U421 ( .A(Packet_In[1]), .Z(n511) );
  N1M1P U422 ( .A(Packet_In[4]), .Z(n517) );
  N1M1P U423 ( .A(Packet_In[13]), .Z(n535) );
  N1M1P U424 ( .A(Packet_In[28]), .Z(n565) );
  N1M1P U425 ( .A(Packet_In[29]), .Z(n567) );
  N1M1P U426 ( .A(Packet_In[26]), .Z(n561) );
  N1M1P U427 ( .A(Packet_In[11]), .Z(n531) );
  N1M1P U428 ( .A(Packet_In[6]), .Z(n521) );
  N1M1P U429 ( .A(Packet_In[22]), .Z(n553) );
  N1M1P U430 ( .A(Packet_In[9]), .Z(n527) );
  N1M1P U431 ( .A(Packet_In[18]), .Z(n545) );
  N1M1P U432 ( .A(Packet_In[23]), .Z(n555) );
  N1M1P U433 ( .A(Packet_In[19]), .Z(n547) );
  N1M1P U434 ( .A(Packet_In[7]), .Z(n523) );
  N1M1P U435 ( .A(Packet_In[10]), .Z(n529) );
  N1M1P U436 ( .A(Packet_In[21]), .Z(n551) );
  N1M1P U437 ( .A(Packet_In[20]), .Z(n549) );
  NR2M1P U438 ( .A(n502), .B(Write_Ack), .Z(n573) );
  NR2M1P U439 ( .A(n392), .B(n573), .Z(n572) );
  AOI22CDNM1P U440 ( .A(n572), .B(n396), .C(n572), .D(n396), .Z(n372) );
  N1M1P U441 ( .A(n573), .Z(n391) );
  AOI22M1P U442 ( .A(Count[0]), .B(n504), .C(n391), .D(n396), .Z(n388) );
  AOI22CDNM1P U443 ( .A(Count[1]), .B(n388), .C(n388), .D(Count[1]), .Z(n371)
         );
  ND2M1P U444 ( .A(Count[1]), .B(Read_Ack), .Z(n387) );
  OAI211M1P U445 ( .A(Count[1]), .B(n504), .C(n388), .D(n387), .Z(n389) );
  AOI22M1P U446 ( .A(n392), .B(n505), .C(Count[2]), .D(n389), .Z(n390) );
  OAI21M1P U447 ( .A(n430), .B(n391), .C(n390), .Z(n370) );
  AOI22CDNM1P U448 ( .A(n383), .B(n571), .C(\Queue[4][31] ), .D(n383), .Z(n369) );
  AOI22CDNM1P U449 ( .A(n383), .B(n509), .C(\Queue[4][0] ), .D(n383), .Z(n368)
         );
  AOI22CDNM1P U450 ( .A(n383), .B(n511), .C(\Queue[4][1] ), .D(n383), .Z(n367)
         );
  AOI22CDNM1P U451 ( .A(n383), .B(n513), .C(\Queue[4][2] ), .D(n383), .Z(n366)
         );
  AOI22CDNM1P U452 ( .A(n383), .B(n515), .C(\Queue[4][3] ), .D(n383), .Z(n365)
         );
  AOI22CDNM1P U453 ( .A(n383), .B(n517), .C(\Queue[4][4] ), .D(n383), .Z(n364)
         );
  AOI22CDNM1P U454 ( .A(n383), .B(n519), .C(\Queue[4][5] ), .D(n383), .Z(n363)
         );
  AOI22CDNM1P U455 ( .A(n383), .B(n521), .C(\Queue[4][6] ), .D(n383), .Z(n362)
         );
  AOI22CDNM1P U456 ( .A(n383), .B(n523), .C(\Queue[4][7] ), .D(n383), .Z(n361)
         );
  AOI22CDNM1P U457 ( .A(n383), .B(n525), .C(\Queue[4][8] ), .D(n383), .Z(n360)
         );
  AOI22CDNM1P U458 ( .A(n383), .B(n527), .C(\Queue[4][9] ), .D(n383), .Z(n359)
         );
  AOI22CDNM1P U459 ( .A(n383), .B(n529), .C(\Queue[4][10] ), .D(n383), .Z(n358) );
  AOI22CDNM1P U460 ( .A(n383), .B(n531), .C(\Queue[4][11] ), .D(n383), .Z(n357) );
  AOI22CDNM1P U461 ( .A(n383), .B(n533), .C(\Queue[4][12] ), .D(n383), .Z(n356) );
  AOI22CDNM1P U462 ( .A(n383), .B(n535), .C(\Queue[4][13] ), .D(n383), .Z(n355) );
  AOI22CDNM1P U463 ( .A(n383), .B(n537), .C(\Queue[4][14] ), .D(n383), .Z(n354) );
  AOI22CDNM1P U464 ( .A(n383), .B(n539), .C(\Queue[4][15] ), .D(n383), .Z(n353) );
  AOI22CDNM1P U465 ( .A(n383), .B(n541), .C(\Queue[4][16] ), .D(n383), .Z(n352) );
  AOI22CDNM1P U466 ( .A(n383), .B(n543), .C(\Queue[4][17] ), .D(n383), .Z(n351) );
  AOI22CDNM1P U467 ( .A(n383), .B(n545), .C(\Queue[4][18] ), .D(n383), .Z(n350) );
  AOI22CDNM1P U468 ( .A(n383), .B(n547), .C(\Queue[4][19] ), .D(n383), .Z(n349) );
  AOI22CDNM1P U469 ( .A(n383), .B(n549), .C(\Queue[4][20] ), .D(n383), .Z(n348) );
  AOI22CDNM1P U470 ( .A(n383), .B(n551), .C(\Queue[4][21] ), .D(n383), .Z(n347) );
  AOI22CDNM1P U471 ( .A(n383), .B(n553), .C(\Queue[4][22] ), .D(n383), .Z(n346) );
  AOI22CDNM1P U472 ( .A(n383), .B(n555), .C(\Queue[4][23] ), .D(n383), .Z(n345) );
  AOI22CDNM1P U473 ( .A(n383), .B(n557), .C(\Queue[4][24] ), .D(n383), .Z(n344) );
  AOI22CDNM1P U474 ( .A(n383), .B(n559), .C(\Queue[4][25] ), .D(n383), .Z(n343) );
  AOI22CDNM1P U475 ( .A(n383), .B(n561), .C(\Queue[4][26] ), .D(n383), .Z(n342) );
  AOI22CDNM1P U476 ( .A(n383), .B(n563), .C(\Queue[4][27] ), .D(n383), .Z(n341) );
  AOI22CDNM1P U477 ( .A(n383), .B(n565), .C(\Queue[4][28] ), .D(n383), .Z(n340) );
  AOI22CDNM1P U478 ( .A(n383), .B(n567), .C(\Queue[4][29] ), .D(n383), .Z(n339) );
  AOI22CDNM1P U479 ( .A(n383), .B(n569), .C(\Queue[4][30] ), .D(n383), .Z(n338) );
  OAI22CDNM1P U480 ( .A(n504), .B(n394), .C(n572), .D(Full), .Z(n337) );
  OA21M1P U481 ( .A(n504), .B(n574), .C(Rst_n), .Z(n397) );
  AOI22M1P U482 ( .A(\Queue[2][0] ), .B(n378), .C(\Queue[1][0] ), .D(n385), 
        .Z(n398) );
  OAI21M1P U483 ( .A(n509), .B(n374), .C(n398), .Z(n336) );
  AOI22M1P U484 ( .A(n378), .B(\Queue[2][1] ), .C(\Queue[1][1] ), .D(n385), 
        .Z(n399) );
  OAI21M1P U485 ( .A(n374), .B(n511), .C(n399), .Z(n335) );
  AOI22M1P U486 ( .A(n378), .B(\Queue[2][2] ), .C(\Queue[1][2] ), .D(n385), 
        .Z(n400) );
  OAI21M1P U487 ( .A(n374), .B(n513), .C(n400), .Z(n334) );
  AOI22M1P U488 ( .A(n378), .B(\Queue[2][3] ), .C(\Queue[1][3] ), .D(n385), 
        .Z(n401) );
  OAI21M1P U489 ( .A(n374), .B(n515), .C(n401), .Z(n333) );
  AOI22M1P U490 ( .A(n378), .B(\Queue[2][4] ), .C(\Queue[1][4] ), .D(n385), 
        .Z(n402) );
  OAI21M1P U491 ( .A(n374), .B(n517), .C(n402), .Z(n332) );
  AOI22M1P U492 ( .A(n378), .B(\Queue[2][5] ), .C(\Queue[1][5] ), .D(n385), 
        .Z(n403) );
  OAI21M1P U493 ( .A(n374), .B(n519), .C(n403), .Z(n331) );
  AOI22M1P U494 ( .A(n378), .B(\Queue[2][6] ), .C(\Queue[1][6] ), .D(n385), 
        .Z(n404) );
  OAI21M1P U495 ( .A(n374), .B(n521), .C(n404), .Z(n330) );
  AOI22M1P U496 ( .A(n378), .B(\Queue[2][7] ), .C(\Queue[1][7] ), .D(n385), 
        .Z(n405) );
  OAI21M1P U497 ( .A(n374), .B(n523), .C(n405), .Z(n329) );
  AOI22M1P U498 ( .A(n378), .B(\Queue[2][8] ), .C(\Queue[1][8] ), .D(n385), 
        .Z(n406) );
  OAI21M1P U499 ( .A(n374), .B(n525), .C(n406), .Z(n328) );
  AOI22M1P U500 ( .A(n378), .B(\Queue[2][9] ), .C(\Queue[1][9] ), .D(n385), 
        .Z(n407) );
  OAI21M1P U501 ( .A(n374), .B(n527), .C(n407), .Z(n327) );
  AOI22M1P U502 ( .A(n378), .B(\Queue[2][10] ), .C(\Queue[1][10] ), .D(n385), 
        .Z(n408) );
  OAI21M1P U503 ( .A(n374), .B(n529), .C(n408), .Z(n326) );
  AOI22M1P U504 ( .A(n378), .B(\Queue[2][11] ), .C(\Queue[1][11] ), .D(n385), 
        .Z(n409) );
  OAI21M1P U505 ( .A(n374), .B(n531), .C(n409), .Z(n325) );
  AOI22M1P U506 ( .A(n378), .B(\Queue[2][12] ), .C(\Queue[1][12] ), .D(n385), 
        .Z(n410) );
  OAI21M1P U507 ( .A(n374), .B(n533), .C(n410), .Z(n324) );
  AOI22M1P U508 ( .A(n378), .B(\Queue[2][13] ), .C(\Queue[1][13] ), .D(n385), 
        .Z(n411) );
  OAI21M1P U509 ( .A(n374), .B(n535), .C(n411), .Z(n323) );
  AOI22M1P U510 ( .A(n378), .B(\Queue[2][14] ), .C(\Queue[1][14] ), .D(n385), 
        .Z(n412) );
  OAI21M1P U511 ( .A(n374), .B(n537), .C(n412), .Z(n322) );
  AOI22M1P U512 ( .A(n378), .B(\Queue[2][15] ), .C(\Queue[1][15] ), .D(n385), 
        .Z(n413) );
  OAI21M1P U513 ( .A(n374), .B(n539), .C(n413), .Z(n321) );
  AOI22M1P U514 ( .A(n378), .B(\Queue[2][16] ), .C(\Queue[1][16] ), .D(n385), 
        .Z(n414) );
  OAI21M1P U515 ( .A(n374), .B(n541), .C(n414), .Z(n320) );
  AOI22M1P U516 ( .A(n378), .B(\Queue[2][17] ), .C(\Queue[1][17] ), .D(n385), 
        .Z(n415) );
  OAI21M1P U517 ( .A(n374), .B(n543), .C(n415), .Z(n319) );
  AOI22M1P U518 ( .A(n378), .B(\Queue[2][18] ), .C(\Queue[1][18] ), .D(n385), 
        .Z(n416) );
  OAI21M1P U519 ( .A(n374), .B(n545), .C(n416), .Z(n318) );
  AOI22M1P U520 ( .A(n378), .B(\Queue[2][19] ), .C(\Queue[1][19] ), .D(n385), 
        .Z(n417) );
  OAI21M1P U521 ( .A(n374), .B(n547), .C(n417), .Z(n317) );
  AOI22M1P U522 ( .A(n378), .B(\Queue[2][20] ), .C(\Queue[1][20] ), .D(n385), 
        .Z(n418) );
  OAI21M1P U523 ( .A(n374), .B(n549), .C(n418), .Z(n316) );
  AOI22M1P U524 ( .A(n378), .B(\Queue[2][21] ), .C(\Queue[1][21] ), .D(n385), 
        .Z(n419) );
  OAI21M1P U525 ( .A(n374), .B(n551), .C(n419), .Z(n315) );
  AOI22M1P U526 ( .A(n378), .B(\Queue[2][22] ), .C(\Queue[1][22] ), .D(n385), 
        .Z(n420) );
  OAI21M1P U527 ( .A(n374), .B(n553), .C(n420), .Z(n314) );
  AOI22M1P U528 ( .A(n378), .B(\Queue[2][23] ), .C(\Queue[1][23] ), .D(n385), 
        .Z(n421) );
  OAI21M1P U529 ( .A(n374), .B(n555), .C(n421), .Z(n313) );
  AOI22M1P U530 ( .A(n378), .B(\Queue[2][24] ), .C(\Queue[1][24] ), .D(n385), 
        .Z(n422) );
  OAI21M1P U531 ( .A(n374), .B(n557), .C(n422), .Z(n312) );
  AOI22M1P U532 ( .A(n378), .B(\Queue[2][25] ), .C(\Queue[1][25] ), .D(n385), 
        .Z(n423) );
  OAI21M1P U533 ( .A(n374), .B(n559), .C(n423), .Z(n311) );
  AOI22M1P U534 ( .A(n378), .B(\Queue[2][26] ), .C(\Queue[1][26] ), .D(n385), 
        .Z(n424) );
  OAI21M1P U535 ( .A(n374), .B(n561), .C(n424), .Z(n310) );
  AOI22M1P U536 ( .A(n378), .B(\Queue[2][27] ), .C(\Queue[1][27] ), .D(n385), 
        .Z(n425) );
  OAI21M1P U537 ( .A(n374), .B(n563), .C(n425), .Z(n309) );
  AOI22M1P U538 ( .A(n378), .B(\Queue[2][28] ), .C(\Queue[1][28] ), .D(n385), 
        .Z(n426) );
  OAI21M1P U539 ( .A(n374), .B(n565), .C(n426), .Z(n308) );
  AOI22M1P U540 ( .A(n378), .B(\Queue[2][29] ), .C(\Queue[1][29] ), .D(n385), 
        .Z(n427) );
  OAI21M1P U541 ( .A(n374), .B(n567), .C(n427), .Z(n307) );
  AOI22M1P U542 ( .A(n378), .B(\Queue[2][30] ), .C(\Queue[1][30] ), .D(n385), 
        .Z(n428) );
  OAI21M1P U543 ( .A(n374), .B(n569), .C(n428), .Z(n306) );
  AOI22M1P U544 ( .A(n378), .B(\Queue[2][31] ), .C(\Queue[1][31] ), .D(n385), 
        .Z(n429) );
  OAI21M1P U545 ( .A(n374), .B(n571), .C(n429), .Z(n305) );
  AOI22M1P U546 ( .A(\Queue[1][0] ), .B(n379), .C(n386), .D(Packet_Out[0]), 
        .Z(n433) );
  OAI21M1P U547 ( .A(n509), .B(n376), .C(n433), .Z(n304) );
  AOI22M1P U548 ( .A(\Queue[1][1] ), .B(n379), .C(n386), .D(Packet_Out[1]), 
        .Z(n434) );
  OAI21M1P U549 ( .A(n511), .B(n376), .C(n434), .Z(n303) );
  AOI22M1P U550 ( .A(\Queue[1][2] ), .B(n379), .C(n386), .D(Packet_Out[2]), 
        .Z(n435) );
  OAI21M1P U551 ( .A(n513), .B(n376), .C(n435), .Z(n302) );
  AOI22M1P U552 ( .A(\Queue[1][3] ), .B(n379), .C(n386), .D(Packet_Out[3]), 
        .Z(n436) );
  OAI21M1P U553 ( .A(n515), .B(n376), .C(n436), .Z(n301) );
  AOI22M1P U554 ( .A(\Queue[1][4] ), .B(n379), .C(n386), .D(Packet_Out[4]), 
        .Z(n437) );
  OAI21M1P U555 ( .A(n517), .B(n376), .C(n437), .Z(n300) );
  AOI22M1P U556 ( .A(\Queue[1][5] ), .B(n379), .C(n386), .D(Packet_Out[5]), 
        .Z(n438) );
  OAI21M1P U557 ( .A(n519), .B(n376), .C(n438), .Z(n299) );
  AOI22M1P U558 ( .A(\Queue[1][6] ), .B(n379), .C(n386), .D(Packet_Out[6]), 
        .Z(n439) );
  OAI21M1P U559 ( .A(n521), .B(n376), .C(n439), .Z(n298) );
  AOI22M1P U560 ( .A(\Queue[1][7] ), .B(n379), .C(n386), .D(Packet_Out[7]), 
        .Z(n440) );
  OAI21M1P U561 ( .A(n523), .B(n376), .C(n440), .Z(n297) );
  AOI22M1P U562 ( .A(\Queue[1][8] ), .B(n379), .C(n464), .D(Packet_Out[8]), 
        .Z(n441) );
  OAI21M1P U563 ( .A(n525), .B(n376), .C(n441), .Z(n296) );
  AOI22M1P U564 ( .A(\Queue[1][9] ), .B(n379), .C(n464), .D(Packet_Out[9]), 
        .Z(n442) );
  OAI21M1P U565 ( .A(n527), .B(n376), .C(n442), .Z(n295) );
  AOI22M1P U566 ( .A(\Queue[1][10] ), .B(n379), .C(n386), .D(Packet_Out[10]), 
        .Z(n443) );
  OAI21M1P U567 ( .A(n529), .B(n376), .C(n443), .Z(n294) );
  AOI22M1P U568 ( .A(\Queue[1][11] ), .B(n379), .C(n386), .D(Packet_Out[11]), 
        .Z(n444) );
  OAI21M1P U569 ( .A(n531), .B(n376), .C(n444), .Z(n293) );
  AOI22M1P U570 ( .A(\Queue[1][12] ), .B(n379), .C(n464), .D(Packet_Out[12]), 
        .Z(n445) );
  OAI21M1P U571 ( .A(n533), .B(n376), .C(n445), .Z(n292) );
  AOI22M1P U572 ( .A(\Queue[1][13] ), .B(n379), .C(n386), .D(Packet_Out[13]), 
        .Z(n446) );
  OAI21M1P U573 ( .A(n535), .B(n376), .C(n446), .Z(n291) );
  AOI22M1P U574 ( .A(\Queue[1][14] ), .B(n379), .C(n464), .D(Packet_Out[14]), 
        .Z(n447) );
  OAI21M1P U575 ( .A(n537), .B(n376), .C(n447), .Z(n290) );
  AOI22M1P U576 ( .A(\Queue[1][15] ), .B(n379), .C(n386), .D(Packet_Out[15]), 
        .Z(n448) );
  OAI21M1P U577 ( .A(n539), .B(n376), .C(n448), .Z(n289) );
  AOI22M1P U578 ( .A(\Queue[1][16] ), .B(n379), .C(n464), .D(Packet_Out[16]), 
        .Z(n449) );
  OAI21M1P U579 ( .A(n541), .B(n376), .C(n449), .Z(n288) );
  AOI22M1P U580 ( .A(\Queue[1][17] ), .B(n379), .C(n464), .D(Packet_Out[17]), 
        .Z(n450) );
  OAI21M1P U581 ( .A(n543), .B(n376), .C(n450), .Z(n287) );
  AOI22M1P U582 ( .A(\Queue[1][18] ), .B(n379), .C(n386), .D(Packet_Out[18]), 
        .Z(n451) );
  OAI21M1P U583 ( .A(n545), .B(n376), .C(n451), .Z(n286) );
  AOI22M1P U584 ( .A(\Queue[1][19] ), .B(n379), .C(n386), .D(Packet_Out[19]), 
        .Z(n452) );
  OAI21M1P U585 ( .A(n547), .B(n376), .C(n452), .Z(n285) );
  AOI22M1P U586 ( .A(\Queue[1][20] ), .B(n379), .C(n464), .D(Packet_Out[20]), 
        .Z(n453) );
  OAI21M1P U587 ( .A(n549), .B(n376), .C(n453), .Z(n284) );
  AOI22M1P U588 ( .A(\Queue[1][21] ), .B(n379), .C(n386), .D(Packet_Out[21]), 
        .Z(n454) );
  OAI21M1P U589 ( .A(n551), .B(n376), .C(n454), .Z(n283) );
  AOI22M1P U590 ( .A(\Queue[1][22] ), .B(n379), .C(n386), .D(Packet_Out[22]), 
        .Z(n455) );
  OAI21M1P U591 ( .A(n553), .B(n376), .C(n455), .Z(n282) );
  AOI22M1P U592 ( .A(\Queue[1][23] ), .B(n379), .C(n464), .D(Packet_Out[23]), 
        .Z(n456) );
  OAI21M1P U593 ( .A(n555), .B(n376), .C(n456), .Z(n281) );
  AOI22M1P U594 ( .A(\Queue[1][24] ), .B(n379), .C(n464), .D(Packet_Out[24]), 
        .Z(n457) );
  OAI21M1P U595 ( .A(n557), .B(n376), .C(n457), .Z(n280) );
  AOI22M1P U596 ( .A(\Queue[1][25] ), .B(n379), .C(n464), .D(Packet_Out[25]), 
        .Z(n458) );
  OAI21M1P U597 ( .A(n559), .B(n376), .C(n458), .Z(n279) );
  AOI22M1P U598 ( .A(\Queue[1][26] ), .B(n379), .C(n386), .D(Packet_Out[26]), 
        .Z(n459) );
  OAI21M1P U599 ( .A(n561), .B(n376), .C(n459), .Z(n278) );
  AOI22M1P U600 ( .A(\Queue[1][27] ), .B(n379), .C(n386), .D(Packet_Out[27]), 
        .Z(n460) );
  OAI21M1P U601 ( .A(n563), .B(n376), .C(n460), .Z(n277) );
  AOI22M1P U602 ( .A(\Queue[1][28] ), .B(n379), .C(n386), .D(Packet_Out[28]), 
        .Z(n461) );
  OAI21M1P U603 ( .A(n565), .B(n376), .C(n461), .Z(n276) );
  AOI22M1P U604 ( .A(\Queue[1][29] ), .B(n379), .C(n386), .D(Packet_Out[29]), 
        .Z(n462) );
  OAI21M1P U605 ( .A(n567), .B(n376), .C(n462), .Z(n275) );
  AOI22M1P U606 ( .A(\Queue[1][30] ), .B(n379), .C(n386), .D(Packet_Out[30]), 
        .Z(n463) );
  OAI21M1P U607 ( .A(n569), .B(n376), .C(n463), .Z(n274) );
  AOI22M1P U608 ( .A(\Queue[1][31] ), .B(n379), .C(n386), .D(Packet_Out[31]), 
        .Z(n465) );
  OAI21M1P U609 ( .A(n571), .B(n376), .C(n465), .Z(n273) );
  OA21M1P U610 ( .A(n504), .B(n468), .C(Rst_n), .Z(n466) );
  ND2M1P U611 ( .A(n467), .B(n502), .Z(n503) );
  AOI22M1P U612 ( .A(\Queue[2][0] ), .B(n375), .C(\Queue[3][0] ), .D(n380), 
        .Z(n469) );
  OAI21M1P U613 ( .A(n509), .B(n373), .C(n469), .Z(n272) );
  AOI22M1P U614 ( .A(\Queue[2][1] ), .B(n375), .C(n380), .D(\Queue[3][1] ), 
        .Z(n470) );
  OAI21M1P U615 ( .A(n511), .B(n373), .C(n470), .Z(n271) );
  AOI22M1P U616 ( .A(\Queue[2][2] ), .B(n375), .C(n380), .D(\Queue[3][2] ), 
        .Z(n471) );
  OAI21M1P U617 ( .A(n513), .B(n373), .C(n471), .Z(n270) );
  AOI22M1P U618 ( .A(\Queue[2][3] ), .B(n375), .C(n380), .D(\Queue[3][3] ), 
        .Z(n472) );
  OAI21M1P U619 ( .A(n515), .B(n373), .C(n472), .Z(n269) );
  AOI22M1P U620 ( .A(\Queue[2][4] ), .B(n375), .C(n380), .D(\Queue[3][4] ), 
        .Z(n473) );
  OAI21M1P U621 ( .A(n517), .B(n373), .C(n473), .Z(n268) );
  AOI22M1P U622 ( .A(\Queue[2][5] ), .B(n375), .C(n380), .D(\Queue[3][5] ), 
        .Z(n474) );
  OAI21M1P U623 ( .A(n519), .B(n373), .C(n474), .Z(n267) );
  AOI22M1P U624 ( .A(\Queue[2][6] ), .B(n375), .C(n380), .D(\Queue[3][6] ), 
        .Z(n475) );
  OAI21M1P U625 ( .A(n521), .B(n373), .C(n475), .Z(n266) );
  AOI22M1P U626 ( .A(\Queue[2][7] ), .B(n375), .C(n380), .D(\Queue[3][7] ), 
        .Z(n476) );
  OAI21M1P U627 ( .A(n523), .B(n373), .C(n476), .Z(n265) );
  AOI22M1P U628 ( .A(\Queue[2][8] ), .B(n375), .C(n380), .D(\Queue[3][8] ), 
        .Z(n477) );
  OAI21M1P U629 ( .A(n525), .B(n373), .C(n477), .Z(n264) );
  AOI22M1P U630 ( .A(\Queue[2][9] ), .B(n375), .C(n380), .D(\Queue[3][9] ), 
        .Z(n478) );
  OAI21M1P U631 ( .A(n527), .B(n373), .C(n478), .Z(n263) );
  AOI22M1P U632 ( .A(\Queue[2][10] ), .B(n375), .C(n380), .D(\Queue[3][10] ), 
        .Z(n479) );
  OAI21M1P U633 ( .A(n529), .B(n373), .C(n479), .Z(n262) );
  AOI22M1P U634 ( .A(\Queue[2][11] ), .B(n375), .C(n380), .D(\Queue[3][11] ), 
        .Z(n480) );
  OAI21M1P U635 ( .A(n531), .B(n373), .C(n480), .Z(n261) );
  AOI22M1P U636 ( .A(\Queue[2][12] ), .B(n375), .C(n380), .D(\Queue[3][12] ), 
        .Z(n481) );
  OAI21M1P U637 ( .A(n533), .B(n373), .C(n481), .Z(n260) );
  AOI22M1P U638 ( .A(\Queue[2][13] ), .B(n375), .C(n380), .D(\Queue[3][13] ), 
        .Z(n482) );
  OAI21M1P U639 ( .A(n535), .B(n373), .C(n482), .Z(n259) );
  AOI22M1P U640 ( .A(\Queue[2][14] ), .B(n375), .C(n380), .D(\Queue[3][14] ), 
        .Z(n483) );
  OAI21M1P U641 ( .A(n537), .B(n373), .C(n483), .Z(n258) );
  AOI22M1P U642 ( .A(\Queue[2][15] ), .B(n375), .C(n380), .D(\Queue[3][15] ), 
        .Z(n484) );
  OAI21M1P U643 ( .A(n539), .B(n373), .C(n484), .Z(n257) );
  AOI22M1P U644 ( .A(\Queue[2][16] ), .B(n375), .C(n380), .D(\Queue[3][16] ), 
        .Z(n485) );
  OAI21M1P U645 ( .A(n541), .B(n373), .C(n485), .Z(n256) );
  AOI22M1P U646 ( .A(\Queue[2][17] ), .B(n375), .C(n380), .D(\Queue[3][17] ), 
        .Z(n486) );
  OAI21M1P U647 ( .A(n543), .B(n373), .C(n486), .Z(n255) );
  AOI22M1P U648 ( .A(\Queue[2][18] ), .B(n375), .C(n380), .D(\Queue[3][18] ), 
        .Z(n487) );
  OAI21M1P U649 ( .A(n545), .B(n373), .C(n487), .Z(n254) );
  AOI22M1P U650 ( .A(\Queue[2][19] ), .B(n375), .C(n380), .D(\Queue[3][19] ), 
        .Z(n488) );
  OAI21M1P U651 ( .A(n547), .B(n373), .C(n488), .Z(n253) );
  AOI22M1P U652 ( .A(\Queue[2][20] ), .B(n375), .C(n380), .D(\Queue[3][20] ), 
        .Z(n489) );
  OAI21M1P U653 ( .A(n549), .B(n373), .C(n489), .Z(n252) );
  AOI22M1P U654 ( .A(\Queue[2][21] ), .B(n375), .C(n380), .D(\Queue[3][21] ), 
        .Z(n490) );
  OAI21M1P U655 ( .A(n551), .B(n373), .C(n490), .Z(n251) );
  AOI22M1P U656 ( .A(\Queue[2][22] ), .B(n375), .C(n380), .D(\Queue[3][22] ), 
        .Z(n491) );
  OAI21M1P U657 ( .A(n553), .B(n373), .C(n491), .Z(n250) );
  AOI22M1P U658 ( .A(\Queue[2][23] ), .B(n375), .C(n380), .D(\Queue[3][23] ), 
        .Z(n492) );
  OAI21M1P U659 ( .A(n555), .B(n373), .C(n492), .Z(n249) );
  AOI22M1P U660 ( .A(\Queue[2][24] ), .B(n375), .C(n380), .D(\Queue[3][24] ), 
        .Z(n493) );
  OAI21M1P U661 ( .A(n557), .B(n373), .C(n493), .Z(n248) );
  AOI22M1P U662 ( .A(\Queue[2][25] ), .B(n375), .C(n380), .D(\Queue[3][25] ), 
        .Z(n494) );
  OAI21M1P U663 ( .A(n559), .B(n373), .C(n494), .Z(n247) );
  AOI22M1P U664 ( .A(\Queue[2][26] ), .B(n375), .C(n380), .D(\Queue[3][26] ), 
        .Z(n495) );
  OAI21M1P U665 ( .A(n561), .B(n373), .C(n495), .Z(n246) );
  AOI22M1P U666 ( .A(\Queue[2][27] ), .B(n375), .C(n380), .D(\Queue[3][27] ), 
        .Z(n496) );
  OAI21M1P U667 ( .A(n563), .B(n373), .C(n496), .Z(n245) );
  AOI22M1P U668 ( .A(\Queue[2][28] ), .B(n375), .C(n380), .D(\Queue[3][28] ), 
        .Z(n497) );
  OAI21M1P U669 ( .A(n565), .B(n373), .C(n497), .Z(n244) );
  AOI22M1P U670 ( .A(\Queue[2][29] ), .B(n375), .C(n380), .D(\Queue[3][29] ), 
        .Z(n498) );
  OAI21M1P U671 ( .A(n567), .B(n373), .C(n498), .Z(n243) );
  AOI22M1P U672 ( .A(\Queue[2][30] ), .B(n375), .C(n380), .D(\Queue[3][30] ), 
        .Z(n499) );
  OAI21M1P U673 ( .A(n569), .B(n373), .C(n499), .Z(n242) );
  AOI22M1P U674 ( .A(\Queue[2][31] ), .B(n375), .C(n380), .D(\Queue[3][31] ), 
        .Z(n500) );
  OAI21M1P U675 ( .A(n571), .B(n373), .C(n500), .Z(n241) );
  OA21M1P U676 ( .A(n504), .B(n505), .C(Rst_n), .Z(n501) );
  AOI22M1P U677 ( .A(\Queue[3][0] ), .B(n382), .C(n381), .D(\Queue[4][0] ), 
        .Z(n508) );
  OAI21M1P U678 ( .A(n509), .B(n377), .C(n508), .Z(n240) );
  AOI22M1P U679 ( .A(\Queue[3][1] ), .B(n382), .C(n381), .D(\Queue[4][1] ), 
        .Z(n510) );
  OAI21M1P U680 ( .A(n511), .B(n377), .C(n510), .Z(n239) );
  AOI22M1P U681 ( .A(\Queue[3][2] ), .B(n382), .C(n381), .D(\Queue[4][2] ), 
        .Z(n512) );
  OAI21M1P U682 ( .A(n513), .B(n377), .C(n512), .Z(n238) );
  AOI22M1P U683 ( .A(\Queue[3][3] ), .B(n382), .C(n381), .D(\Queue[4][3] ), 
        .Z(n514) );
  OAI21M1P U684 ( .A(n515), .B(n377), .C(n514), .Z(n237) );
  AOI22M1P U685 ( .A(\Queue[3][4] ), .B(n382), .C(n381), .D(\Queue[4][4] ), 
        .Z(n516) );
  OAI21M1P U686 ( .A(n517), .B(n377), .C(n516), .Z(n236) );
  AOI22M1P U687 ( .A(\Queue[3][5] ), .B(n382), .C(n381), .D(\Queue[4][5] ), 
        .Z(n518) );
  OAI21M1P U688 ( .A(n519), .B(n377), .C(n518), .Z(n235) );
  AOI22M1P U689 ( .A(\Queue[3][6] ), .B(n382), .C(n381), .D(\Queue[4][6] ), 
        .Z(n520) );
  OAI21M1P U690 ( .A(n521), .B(n377), .C(n520), .Z(n234) );
  AOI22M1P U691 ( .A(\Queue[3][7] ), .B(n382), .C(n381), .D(\Queue[4][7] ), 
        .Z(n522) );
  OAI21M1P U692 ( .A(n523), .B(n377), .C(n522), .Z(n233) );
  AOI22M1P U693 ( .A(\Queue[3][8] ), .B(n382), .C(n381), .D(\Queue[4][8] ), 
        .Z(n524) );
  OAI21M1P U694 ( .A(n525), .B(n377), .C(n524), .Z(n232) );
  AOI22M1P U695 ( .A(\Queue[3][9] ), .B(n382), .C(n381), .D(\Queue[4][9] ), 
        .Z(n526) );
  OAI21M1P U696 ( .A(n527), .B(n377), .C(n526), .Z(n231) );
  AOI22M1P U697 ( .A(\Queue[3][10] ), .B(n382), .C(n381), .D(\Queue[4][10] ), 
        .Z(n528) );
  OAI21M1P U698 ( .A(n529), .B(n377), .C(n528), .Z(n230) );
  AOI22M1P U699 ( .A(\Queue[3][11] ), .B(n382), .C(n381), .D(\Queue[4][11] ), 
        .Z(n530) );
  OAI21M1P U700 ( .A(n531), .B(n377), .C(n530), .Z(n229) );
  AOI22M1P U701 ( .A(\Queue[3][12] ), .B(n382), .C(n381), .D(\Queue[4][12] ), 
        .Z(n532) );
  OAI21M1P U702 ( .A(n533), .B(n377), .C(n532), .Z(n228) );
  AOI22M1P U703 ( .A(\Queue[3][13] ), .B(n382), .C(n381), .D(\Queue[4][13] ), 
        .Z(n534) );
  OAI21M1P U704 ( .A(n535), .B(n377), .C(n534), .Z(n227) );
  AOI22M1P U705 ( .A(\Queue[3][14] ), .B(n382), .C(n381), .D(\Queue[4][14] ), 
        .Z(n536) );
  OAI21M1P U706 ( .A(n537), .B(n377), .C(n536), .Z(n226) );
  AOI22M1P U707 ( .A(\Queue[3][15] ), .B(n382), .C(n381), .D(\Queue[4][15] ), 
        .Z(n538) );
  OAI21M1P U708 ( .A(n539), .B(n377), .C(n538), .Z(n225) );
  AOI22M1P U709 ( .A(\Queue[3][16] ), .B(n382), .C(n381), .D(\Queue[4][16] ), 
        .Z(n540) );
  OAI21M1P U710 ( .A(n541), .B(n377), .C(n540), .Z(n224) );
  AOI22M1P U711 ( .A(\Queue[3][17] ), .B(n382), .C(n381), .D(\Queue[4][17] ), 
        .Z(n542) );
  OAI21M1P U712 ( .A(n543), .B(n377), .C(n542), .Z(n223) );
  AOI22M1P U713 ( .A(\Queue[3][18] ), .B(n382), .C(n381), .D(\Queue[4][18] ), 
        .Z(n544) );
  OAI21M1P U714 ( .A(n545), .B(n377), .C(n544), .Z(n222) );
  AOI22M1P U715 ( .A(\Queue[3][19] ), .B(n382), .C(n381), .D(\Queue[4][19] ), 
        .Z(n546) );
  OAI21M1P U716 ( .A(n547), .B(n377), .C(n546), .Z(n221) );
  AOI22M1P U717 ( .A(\Queue[3][20] ), .B(n382), .C(n381), .D(\Queue[4][20] ), 
        .Z(n548) );
  OAI21M1P U718 ( .A(n549), .B(n377), .C(n548), .Z(n220) );
  AOI22M1P U719 ( .A(\Queue[3][21] ), .B(n382), .C(n381), .D(\Queue[4][21] ), 
        .Z(n550) );
  OAI21M1P U720 ( .A(n551), .B(n377), .C(n550), .Z(n219) );
  AOI22M1P U721 ( .A(\Queue[3][22] ), .B(n382), .C(n381), .D(\Queue[4][22] ), 
        .Z(n552) );
  OAI21M1P U722 ( .A(n553), .B(n377), .C(n552), .Z(n218) );
  AOI22M1P U723 ( .A(\Queue[3][23] ), .B(n382), .C(n381), .D(\Queue[4][23] ), 
        .Z(n554) );
  OAI21M1P U724 ( .A(n555), .B(n377), .C(n554), .Z(n217) );
  AOI22M1P U725 ( .A(\Queue[3][24] ), .B(n382), .C(n381), .D(\Queue[4][24] ), 
        .Z(n556) );
  OAI21M1P U726 ( .A(n557), .B(n377), .C(n556), .Z(n216) );
  AOI22M1P U727 ( .A(\Queue[3][25] ), .B(n382), .C(n381), .D(\Queue[4][25] ), 
        .Z(n558) );
  OAI21M1P U728 ( .A(n559), .B(n377), .C(n558), .Z(n215) );
  AOI22M1P U729 ( .A(\Queue[3][26] ), .B(n382), .C(n381), .D(\Queue[4][26] ), 
        .Z(n560) );
  OAI21M1P U730 ( .A(n561), .B(n377), .C(n560), .Z(n214) );
  AOI22M1P U731 ( .A(\Queue[3][27] ), .B(n382), .C(n381), .D(\Queue[4][27] ), 
        .Z(n562) );
  OAI21M1P U732 ( .A(n563), .B(n377), .C(n562), .Z(n213) );
  AOI22M1P U733 ( .A(\Queue[3][28] ), .B(n382), .C(n381), .D(\Queue[4][28] ), 
        .Z(n564) );
  OAI21M1P U734 ( .A(n565), .B(n377), .C(n564), .Z(n212) );
  AOI22M1P U735 ( .A(\Queue[3][29] ), .B(n382), .C(n381), .D(\Queue[4][29] ), 
        .Z(n566) );
  OAI21M1P U736 ( .A(n567), .B(n377), .C(n566), .Z(n211) );
  AOI22M1P U737 ( .A(\Queue[3][30] ), .B(n382), .C(n381), .D(\Queue[4][30] ), 
        .Z(n568) );
  OAI21M1P U738 ( .A(n569), .B(n377), .C(n568), .Z(n210) );
  AOI22M1P U739 ( .A(\Queue[3][31] ), .B(n382), .C(n381), .D(\Queue[4][31] ), 
        .Z(n570) );
  OAI21M1P U740 ( .A(n571), .B(n377), .C(n570), .Z(n209) );
  N1M1P U741 ( .A(n2), .Z(Empty) );
  AOI22M1P U742 ( .A(n574), .B(n573), .C(n572), .D(Empty), .Z(n1) );
endmodule

