library verilog;
use verilog.vl_types.all;
entity prime_detector_behavioral_structural_tb is
end prime_detector_behavioral_structural_tb;
