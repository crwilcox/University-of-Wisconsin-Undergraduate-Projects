library verilog;
use verilog.vl_types.all;
entity ud_counter_tb is
end ud_counter_tb;
