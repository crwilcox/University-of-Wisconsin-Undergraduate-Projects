library verilog;
use verilog.vl_types.all;
entity p2c_tb is
end p2c_tb;
