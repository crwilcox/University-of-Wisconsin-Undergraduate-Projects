library verilog;
use verilog.vl_types.all;
entity p2_2bit_adder is
end p2_2bit_adder;
