
module tx_synth ( Clk_s, Rst_n, TxData_Valid, TxData, Error_Ack, Rx_Ready, Rx_Error, 
        Tx_Ready, Tx_Error, S_Data );
  input [31:0] TxData;
  input Clk_s, Rst_n, TxData_Valid, Error_Ack, Rx_Ready, Rx_Error;
  output Tx_Ready, Tx_Error, S_Data;
  wire   Tx_Error_Next, N77, N146, N186, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n23, n24, n25, n26, n27, n28, n93,
         n157, n162, N127, N129, N130, N131, N100, N102, N101, N103, N104,
         N105, N106, N107, N108, N109, N110, N119, N120, N121, N122, N125,
         N112, N111, N113, N114, N115, N116, N117, N118, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344;
  wire   [32:0] transmissionPacket;
  wire   [5:0] bitCount;

  FD2QM1P Tx_Error_reg ( .D(Tx_Error_Next), .CP(Clk_s), .CD(Rst_n), .Q(
        Tx_Error) );
  FDN2QM1P Tx_Error_Next_reg ( .D(N77), .CPN(Clk_s), .CD(Rst_n), .Q(
        Tx_Error_Next) );
  FD4QM1P zeroPatternDetected_reg ( .D(n14), .CP(Clk_s), .SD(Rst_n), .Q(n15)
         );
  FD4QM1P DataTxInProg_reg ( .D(n12), .CP(Clk_s), .SD(Rst_n), .Q(n13) );
  FD4QM1P Tx_Ready_reg ( .D(n162), .CP(Clk_s), .SD(Rst_n), .Q(Tx_Ready) );
  FD2QM1P \transmissionPacket_reg[0]  ( .D(n157), .CP(Clk_s), .CD(Rst_n), .Q(
        transmissionPacket[0]) );
  FD2LQM1P \transmissionPacket_reg[1]  ( .D(TxData[0]), .LD(n16), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[1]) );
  FD2LQM1P \transmissionPacket_reg[2]  ( .D(TxData[1]), .LD(n16), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[2]) );
  FD2LQM1P \transmissionPacket_reg[3]  ( .D(TxData[2]), .LD(n16), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[3]) );
  FD2LQM1P \transmissionPacket_reg[4]  ( .D(TxData[3]), .LD(n16), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[4]) );
  FD2LQM1P \transmissionPacket_reg[5]  ( .D(TxData[4]), .LD(n16), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[5]) );
  FD2LQM1P \transmissionPacket_reg[6]  ( .D(TxData[5]), .LD(n16), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[6]) );
  FD2LQM1P \transmissionPacket_reg[7]  ( .D(TxData[6]), .LD(n16), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[7]) );
  FD2LQM1P \transmissionPacket_reg[8]  ( .D(TxData[7]), .LD(n16), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[8]) );
  FD2LQM1P \transmissionPacket_reg[9]  ( .D(TxData[8]), .LD(n16), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[9]) );
  FD2LQM1P \transmissionPacket_reg[10]  ( .D(TxData[9]), .LD(n16), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[10]) );
  FD2LQM1P \transmissionPacket_reg[11]  ( .D(TxData[10]), .LD(n16), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[11]) );
  FD2LQM1P \transmissionPacket_reg[12]  ( .D(TxData[11]), .LD(n16), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[12]) );
  FD2LQM1P \transmissionPacket_reg[13]  ( .D(TxData[12]), .LD(n16), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[13]) );
  FD2LQM1P \transmissionPacket_reg[14]  ( .D(TxData[13]), .LD(n16), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[14]) );
  FD2LQM1P \transmissionPacket_reg[15]  ( .D(TxData[14]), .LD(n16), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[15]) );
  FD2LQM1P \transmissionPacket_reg[16]  ( .D(TxData[15]), .LD(n16), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[16]) );
  FD2LQM1P \transmissionPacket_reg[17]  ( .D(TxData[16]), .LD(n16), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[17]) );
  FD2LQM1P \transmissionPacket_reg[18]  ( .D(TxData[17]), .LD(n16), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[18]) );
  FD2LQM1P \transmissionPacket_reg[19]  ( .D(TxData[18]), .LD(n16), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[19]) );
  FD2LQM1P \transmissionPacket_reg[20]  ( .D(TxData[19]), .LD(n16), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[20]) );
  FD2LQM1P \transmissionPacket_reg[21]  ( .D(TxData[20]), .LD(n16), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[21]) );
  FD2LQM1P \transmissionPacket_reg[22]  ( .D(TxData[21]), .LD(n16), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[22]) );
  FD2LQM1P \transmissionPacket_reg[23]  ( .D(TxData[22]), .LD(n16), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[23]) );
  FD2LQM1P \transmissionPacket_reg[24]  ( .D(TxData[23]), .LD(n16), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[24]) );
  FD2LQM1P \transmissionPacket_reg[25]  ( .D(TxData[24]), .LD(n16), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[25]) );
  FD2LQM1P \transmissionPacket_reg[26]  ( .D(TxData[25]), .LD(n16), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[26]) );
  FD2LQM1P \transmissionPacket_reg[27]  ( .D(TxData[26]), .LD(n16), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[27]) );
  FD2LQM1P \transmissionPacket_reg[28]  ( .D(TxData[27]), .LD(n16), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[28]) );
  FD2LQM1P \transmissionPacket_reg[29]  ( .D(TxData[28]), .LD(n16), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[29]) );
  FD2LQM1P \transmissionPacket_reg[30]  ( .D(TxData[29]), .LD(n16), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[30]) );
  FD2LQM1P \transmissionPacket_reg[31]  ( .D(TxData[30]), .LD(n16), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[31]) );
  FD2LQM1P \transmissionPacket_reg[32]  ( .D(TxData[31]), .LD(n16), .CP(Clk_s), 
        .CD(Rst_n), .Q(transmissionPacket[32]) );
  FD4QM1P \startSequenceCount_reg[1]  ( .D(n10), .CP(Clk_s), .SD(Rst_n), .Q(
        n11) );
  FD4QM1P \startSequenceCount_reg[2]  ( .D(n8), .CP(Clk_s), .SD(Rst_n), .Q(n9)
         );
  FD4QM1P \startSequenceCount_reg[0]  ( .D(n6), .CP(Clk_s), .SD(Rst_n), .Q(n7)
         );
  FD4QM1P startSequence_reg ( .D(n93), .CP(Clk_s), .SD(Rst_n), .Q(n5) );
  FD4QM1P \zeroCount_reg[0]  ( .D(n3), .CP(Clk_s), .SD(Rst_n), .Q(n4) );
  FD4QM1P \zeroCount_reg[1]  ( .D(n1), .CP(Clk_s), .SD(Rst_n), .Q(n2) );
  FD4QM1P S_Data_reg ( .D(N146), .CP(Clk_s), .SD(Rst_n), .Q(S_Data) );
  FD2QM8P \bitCount_reg[0]  ( .D(n23), .CP(Clk_s), .CD(Rst_n), .Q(bitCount[0])
         );
  FD2QM8P \bitCount_reg[1]  ( .D(n24), .CP(Clk_s), .CD(Rst_n), .Q(bitCount[1])
         );
  FD2QM8P \bitCount_reg[5]  ( .D(n28), .CP(Clk_s), .CD(Rst_n), .Q(bitCount[5])
         );
  FD2QM8P \bitCount_reg[2]  ( .D(n25), .CP(Clk_s), .CD(Rst_n), .Q(bitCount[2])
         );
  FD2QM8P \bitCount_reg[3]  ( .D(n26), .CP(Clk_s), .CD(Rst_n), .Q(bitCount[3])
         );
  FD2QM8P \bitCount_reg[4]  ( .D(n27), .CP(Clk_s), .CD(Rst_n), .Q(bitCount[4])
         );
  NR2BNM8P U170 ( .B(bitCount[4]), .A(bitCount[5]), .Z(n276) );
  N1M1P U171 ( .A(bitCount[3]), .Z(n176) );
  NR2M2P U172 ( .A(n229), .B(n230), .Z(n208) );
  NR2M1P U173 ( .A(n280), .B(n177), .Z(n165) );
  NR2M1P U174 ( .A(n265), .B(n282), .Z(n166) );
  AOI22M1P U175 ( .A(transmissionPacket[6]), .B(n165), .C(
        transmissionPacket[4]), .D(n166), .Z(n178) );
  NR2M1P U176 ( .A(n282), .B(n177), .Z(n167) );
  NR2M1P U177 ( .A(n275), .B(n270), .Z(n168) );
  AOI22M1P U178 ( .A(transmissionPacket[8]), .B(n167), .C(
        transmissionPacket[9]), .D(n168), .Z(n179) );
  ND2BNM2P U179 ( .B(n273), .A(n329), .Z(n271) );
  N1M1P U180 ( .A(n270), .Z(n169) );
  N1M1P U181 ( .A(n283), .Z(n170) );
  N1M1P U182 ( .A(n280), .Z(n171) );
  AOI222M1P U183 ( .A(n169), .B(transmissionPacket[5]), .C(n170), .D(
        transmissionPacket[7]), .E(n171), .F(transmissionPacket[6]), .Z(n244)
         );
  OA21M1P U184 ( .A(n331), .B(bitCount[1]), .C(n330), .Z(n172) );
  ND3M1P U185 ( .A(n333), .B(bitCount[0]), .C(bitCount[1]), .Z(n173) );
  AOI22M1P U186 ( .A(bitCount[2]), .B(n172), .C(n327), .D(n173), .Z(n25) );
  AND2M4P U187 ( .A(Tx_Ready), .B(TxData_Valid), .Z(n16) );
  N1M6P U188 ( .A(bitCount[0]), .Z(n273) );
  NR2FM1P U189 ( .A(n340), .B(n4), .Z(n344) );
  ND2BNM2P U190 ( .B(n340), .A(n4), .Z(n341) );
  NR2M2P U191 ( .A(n212), .B(n213), .Z(n211) );
  ND3M3P U192 ( .A(bitCount[2]), .B(n276), .C(n285), .Z(n275) );
  N1M8P U193 ( .A(n331), .Z(n333) );
  ND4M8P U194 ( .A(n15), .B(n5), .C(n338), .D(n286), .Z(n331) );
  NR2M2P U195 ( .A(n224), .B(n225), .Z(n209) );
  OAI22M2P U196 ( .A(n283), .B(n236), .C(n282), .D(n237), .Z(n234) );
  AND2M2P U197 ( .A(n319), .B(n320), .Z(n268) );
  ND3M2P U198 ( .A(n268), .B(bitCount[2]), .C(bitCount[3]), .Z(n263) );
  ND2I1M8P U199 ( .A(n268), .B(n175), .Z(n272) );
  NR2FM1P U200 ( .A(n206), .B(n207), .Z(n205) );
  ND4FM2P U201 ( .A(n208), .B(n209), .C(n210), .D(n211), .Z(n207) );
  ND2M8P U202 ( .A(bitCount[1]), .B(n273), .Z(n280) );
  ND4DNFM4P U203 ( .D(bitCount[3]), .A(n329), .B(n327), .C(n320), .Z(n289) );
  NR3M2P U204 ( .A(n199), .B(n198), .C(n197), .Z(n201) );
  ND4FM2P U205 ( .A(n188), .B(n187), .C(n186), .D(n185), .Z(n197) );
  NR2FM2P U206 ( .A(bitCount[5]), .B(bitCount[4]), .Z(n279) );
  ND2M8P U207 ( .A(bitCount[1]), .B(bitCount[0]), .Z(n270) );
  ND2BNM8P U208 ( .B(bitCount[1]), .A(n273), .Z(n282) );
  ND2FM3P U209 ( .A(n277), .B(n276), .Z(n264) );
  NR2M3P U210 ( .A(bitCount[2]), .B(bitCount[3]), .Z(n277) );
  ND4DNFM4P U211 ( .D(n202), .A(n205), .B(n204), .C(n203), .Z(n340) );
  ND2BNM3P U212 ( .B(bitCount[1]), .A(bitCount[0]), .Z(n283) );
  NR2FM1P U213 ( .A(n218), .B(n219), .Z(n210) );
  N1M2P U214 ( .A(bitCount[4]), .Z(n320) );
  N1M2P U215 ( .A(bitCount[2]), .Z(n327) );
  N1M1P U216 ( .A(n13), .Z(n338) );
  N1M2P U217 ( .A(bitCount[1]), .Z(n329) );
  AOI22M1P U218 ( .A(n262), .B(n343), .C(n344), .D(n2), .Z(n1) );
  ND2M1P U219 ( .A(n341), .B(n342), .Z(n262) );
  OAI211M1P U220 ( .A(n201), .B(n331), .C(n15), .D(n200), .Z(N146) );
  AOI21M1P U221 ( .A(N125), .B(transmissionPacket[7]), .C(n180), .Z(n185) );
  AND4M1P U222 ( .A(n184), .B(n183), .C(n182), .D(n181), .Z(n188) );
  OA21M1P U223 ( .A(n4), .B(n342), .C(n341), .Z(n3) );
  ND2M1P U224 ( .A(N186), .B(transmissionPacket[0]), .Z(n203) );
  ND2M1P U225 ( .A(bitCount[5]), .B(n277), .Z(n266) );
  ND2M1P U226 ( .A(n276), .B(n175), .Z(n177) );
  NR2M1P U227 ( .A(n176), .B(bitCount[2]), .Z(n175) );
  ND2BNM1P U228 ( .B(n282), .A(transmissionPacket[8]), .Z(n245) );
  AOI21M1P U229 ( .A(n214), .B(n215), .C(n284), .Z(n213) );
  ND2BNM1P U230 ( .B(n283), .A(transmissionPacket[23]), .Z(n215) );
  ND2BNM1P U231 ( .B(n282), .A(transmissionPacket[24]), .Z(n214) );
  AOI21M1P U232 ( .A(n216), .B(n217), .C(n274), .Z(n212) );
  ND2BNM1P U233 ( .B(n280), .A(transmissionPacket[18]), .Z(n217) );
  ND2BNM1P U234 ( .B(n283), .A(transmissionPacket[19]), .Z(n216) );
  AOI21M1P U235 ( .A(n220), .B(n221), .C(n275), .Z(n219) );
  ND2BNM1P U236 ( .B(n283), .A(transmissionPacket[11]), .Z(n221) );
  ND2BNM1P U237 ( .B(n270), .A(transmissionPacket[9]), .Z(n220) );
  OAI22M1P U238 ( .A(n275), .B(n222), .C(n278), .D(n223), .Z(n218) );
  ND2BNM1P U239 ( .B(n270), .A(transmissionPacket[29]), .Z(n223) );
  ND2BNM1P U240 ( .B(n282), .A(transmissionPacket[12]), .Z(n222) );
  OAI22M1P U241 ( .A(n274), .B(n226), .C(n278), .D(n227), .Z(n225) );
  ND2BNM1P U242 ( .B(n283), .A(transmissionPacket[31]), .Z(n227) );
  ND2BNM1P U243 ( .B(n270), .A(transmissionPacket[17]), .Z(n226) );
  NR2M1P U244 ( .A(n264), .B(n228), .Z(n224) );
  ND2BNM1P U245 ( .B(n270), .A(transmissionPacket[13]), .Z(n228) );
  AOI21M1P U246 ( .A(n231), .B(n232), .C(n278), .Z(n230) );
  ND2M1P U247 ( .A(n279), .B(n277), .Z(n278) );
  ND2BNM1P U248 ( .B(n280), .A(transmissionPacket[30]), .Z(n232) );
  ND2BNM1P U249 ( .B(n282), .A(transmissionPacket[32]), .Z(n231) );
  NR2M1P U250 ( .A(n264), .B(n233), .Z(n229) );
  NR2M1P U251 ( .A(n234), .B(n235), .Z(n233) );
  NR2BNM1P U252 ( .B(transmissionPacket[14]), .A(n280), .Z(n235) );
  N1M1P U253 ( .A(transmissionPacket[16]), .Z(n237) );
  N1M1P U254 ( .A(transmissionPacket[15]), .Z(n236) );
  AOI21M1P U255 ( .A(n238), .B(n239), .C(n265), .Z(n206) );
  ND2M1P U256 ( .A(n276), .B(n174), .Z(n265) );
  AND2M1P U257 ( .A(bitCount[2]), .B(bitCount[3]), .Z(n174) );
  ND2BNM1P U258 ( .B(n282), .A(transmissionPacket[4]), .Z(n239) );
  NR2M1P U259 ( .A(n240), .B(n241), .Z(n238) );
  NR2BNM1P U260 ( .B(transmissionPacket[2]), .A(n280), .Z(n241) );
  OAI22M1P U261 ( .A(n283), .B(n242), .C(n270), .D(n243), .Z(n240) );
  N1M1P U262 ( .A(transmissionPacket[1]), .Z(n243) );
  N1M1P U263 ( .A(transmissionPacket[3]), .Z(n242) );
  ND2M1P U264 ( .A(n246), .B(n247), .Z(n202) );
  NR3M1P U265 ( .A(n248), .B(n249), .C(n250), .Z(n247) );
  OAI21M1P U266 ( .A(n275), .B(n251), .C(n252), .Z(n250) );
  AND3M1P U267 ( .A(n338), .B(n5), .C(n15), .Z(n252) );
  ND2BNM1P U268 ( .B(n280), .A(transmissionPacket[10]), .Z(n251) );
  NR2M1P U269 ( .A(n281), .B(n253), .Z(n249) );
  ND2BNM1P U270 ( .B(n282), .A(transmissionPacket[28]), .Z(n253) );
  AOI21M1P U271 ( .A(n254), .B(n255), .C(n281), .Z(n248) );
  ND2BNM1P U272 ( .B(n280), .A(transmissionPacket[26]), .Z(n255) );
  ND2BNM1P U273 ( .B(n283), .A(transmissionPacket[27]), .Z(n254) );
  NR2M1P U274 ( .A(n256), .B(n257), .Z(n246) );
  OAI22M1P U275 ( .A(n281), .B(n258), .C(n284), .D(n259), .Z(n257) );
  ND2BNM1P U276 ( .B(n270), .A(transmissionPacket[21]), .Z(n259) );
  ND2BNM1P U277 ( .B(n270), .A(transmissionPacket[25]), .Z(n258) );
  ND3M1P U278 ( .A(bitCount[2]), .B(n279), .C(n285), .Z(n281) );
  N1M1P U279 ( .A(bitCount[3]), .Z(n285) );
  OAI22M1P U280 ( .A(n284), .B(n260), .C(n274), .D(n261), .Z(n256) );
  ND2BNM1P U281 ( .B(n282), .A(transmissionPacket[20]), .Z(n261) );
  ND3M1P U282 ( .A(n279), .B(bitCount[2]), .C(bitCount[3]), .Z(n274) );
  ND2BNM1P U283 ( .B(n280), .A(transmissionPacket[22]), .Z(n260) );
  ND3M1P U284 ( .A(n279), .B(bitCount[3]), .C(n327), .Z(n284) );
  N1M1P U285 ( .A(bitCount[5]), .Z(n319) );
  OAI21M1P U286 ( .A(n323), .B(n331), .C(n15), .Z(n325) );
  NR2M1P U287 ( .A(bitCount[3]), .B(n331), .Z(n324) );
  OAI22M1P U288 ( .A(n330), .B(n329), .C(n273), .D(n328), .Z(n24) );
  NR2M1P U289 ( .A(n271), .B(n177), .Z(N125) );
  NR2M1P U290 ( .A(n270), .B(n177), .Z(N127) );
  AO21M1P U291 ( .A(n244), .B(n245), .C(n177), .Z(n204) );
  NR2M1P U292 ( .A(n280), .B(n264), .Z(N118) );
  NR2M1P U293 ( .A(n271), .B(n264), .Z(N117) );
  NR2M1P U294 ( .A(n282), .B(n264), .Z(N116) );
  NR2M1P U295 ( .A(n270), .B(n263), .Z(N115) );
  NR2M1P U296 ( .A(n280), .B(n263), .Z(N114) );
  NR2M1P U297 ( .A(n263), .B(n271), .Z(N113) );
  NR2M1P U298 ( .A(n272), .B(n270), .Z(N111) );
  NR2M1P U299 ( .A(n282), .B(n263), .Z(N112) );
  ND2M1P U300 ( .A(n179), .B(n178), .Z(n180) );
  NR2M1P U301 ( .A(n280), .B(n275), .Z(N122) );
  NR2M1P U302 ( .A(n271), .B(n275), .Z(N121) );
  NR2M1P U303 ( .A(n282), .B(n275), .Z(N120) );
  NR2M1P U304 ( .A(n270), .B(n264), .Z(N119) );
  AOI22M1P U305 ( .A(transmissionPacket[15]), .B(N117), .C(
        transmissionPacket[14]), .D(N118), .Z(n181) );
  AOI22M1P U306 ( .A(transmissionPacket[17]), .B(N115), .C(
        transmissionPacket[16]), .D(N116), .Z(n182) );
  AOI22M1P U307 ( .A(transmissionPacket[19]), .B(N113), .C(
        transmissionPacket[18]), .D(N114), .Z(n183) );
  AOI22M1P U308 ( .A(transmissionPacket[20]), .B(N112), .C(
        transmissionPacket[21]), .D(N111), .Z(n184) );
  NR2M1P U309 ( .A(n272), .B(n280), .Z(N110) );
  NR2M1P U310 ( .A(n272), .B(n271), .Z(N109) );
  NR2M1P U311 ( .A(n282), .B(n272), .Z(N108) );
  NR2M1P U312 ( .A(n270), .B(n269), .Z(N107) );
  NR2M1P U313 ( .A(n280), .B(n269), .Z(N106) );
  NR2M1P U314 ( .A(n271), .B(n269), .Z(N105) );
  NR2M1P U315 ( .A(n282), .B(n269), .Z(N104) );
  NR2M1P U316 ( .A(n267), .B(n270), .Z(N103) );
  NR2M1P U317 ( .A(n267), .B(n271), .Z(N101) );
  NR2M1P U318 ( .A(n267), .B(n280), .Z(N102) );
  NR2M1P U319 ( .A(n282), .B(n267), .Z(N100) );
  NR2M1P U320 ( .A(n270), .B(n265), .Z(N131) );
  NR2M1P U321 ( .A(n280), .B(n265), .Z(N130) );
  NR2M1P U322 ( .A(n271), .B(n265), .Z(N129) );
  AOI22M1P U323 ( .A(transmissionPacket[11]), .B(N121), .C(
        transmissionPacket[10]), .D(N122), .Z(n186) );
  AOI22M1P U324 ( .A(transmissionPacket[13]), .B(N119), .C(
        transmissionPacket[12]), .D(N120), .Z(n187) );
  AOI22M1P U325 ( .A(transmissionPacket[23]), .B(N109), .C(
        transmissionPacket[22]), .D(N110), .Z(n189) );
  AOI22M1P U326 ( .A(transmissionPacket[25]), .B(N107), .C(
        transmissionPacket[24]), .D(N108), .Z(n190) );
  AOI22M1P U327 ( .A(transmissionPacket[27]), .B(N105), .C(
        transmissionPacket[26]), .D(N106), .Z(n191) );
  AOI22M1P U328 ( .A(transmissionPacket[29]), .B(N103), .C(
        transmissionPacket[28]), .D(N104), .Z(n192) );
  AOI22M1P U329 ( .A(transmissionPacket[30]), .B(N102), .C(
        transmissionPacket[31]), .D(N101), .Z(n193) );
  AOI22M1P U330 ( .A(transmissionPacket[32]), .B(N100), .C(
        transmissionPacket[0]), .D(N186), .Z(n194) );
  AOI22M1P U331 ( .A(transmissionPacket[2]), .B(N130), .C(
        transmissionPacket[1]), .D(N131), .Z(n195) );
  AOI22M1P U332 ( .A(transmissionPacket[5]), .B(N127), .C(
        transmissionPacket[3]), .D(N129), .Z(n196) );
  ND4M1P U333 ( .A(n192), .B(n191), .C(n190), .D(n189), .Z(n198) );
  ND4M1P U334 ( .A(n196), .B(n195), .C(n194), .D(n193), .Z(n199) );
  AO21CNM1P U335 ( .A(n338), .B(n286), .C(n5), .Z(n200) );
  ND2M1P U336 ( .A(n268), .B(n277), .Z(n267) );
  ND3M1P U337 ( .A(bitCount[2]), .B(n268), .C(n285), .Z(n269) );
  NR3M1P U338 ( .A(bitCount[4]), .B(n282), .C(n266), .Z(N186) );
  OAI21M1P U339 ( .A(bitCount[0]), .B(n289), .C(bitCount[5]), .Z(n286) );
  N1M1P U340 ( .A(Error_Ack), .Z(n287) );
  AO21M1P U341 ( .A(Tx_Error), .B(n287), .C(Rx_Error), .Z(N77) );
  N1M1P U342 ( .A(Tx_Ready), .Z(n335) );
  AO21M1P U343 ( .A(n7), .B(n11), .C(n9), .Z(n288) );
  ND3M1P U344 ( .A(Rx_Ready), .B(n335), .C(n288), .Z(n93) );
  OR3M1P U345 ( .A(n289), .B(n319), .C(n273), .Z(n290) );
  AOI21M1P U346 ( .A(n335), .B(n290), .C(TxData_Valid), .Z(n162) );
  N1M1P U347 ( .A(transmissionPacket[0]), .Z(n318) );
  AOI22CDNM1P U348 ( .A(TxData[30]), .B(TxData[31]), .C(TxData[31]), .D(
        TxData[30]), .Z(n309) );
  AOI22CDNM1P U349 ( .A(TxData[24]), .B(TxData[25]), .C(TxData[25]), .D(
        TxData[24]), .Z(n294) );
  AOI22CDNM1P U350 ( .A(TxData[26]), .B(TxData[27]), .C(TxData[27]), .D(
        TxData[26]), .Z(n293) );
  N1M1P U351 ( .A(TxData[28]), .Z(n291) );
  AOI22CDNM1P U352 ( .A(TxData[29]), .B(n291), .C(n291), .D(TxData[29]), .Z(
        n292) );
  EN3M1P U353 ( .A(n294), .B(n293), .C(n292), .Z(n308) );
  AOI22CDNM1P U354 ( .A(TxData[6]), .B(TxData[7]), .C(TxData[7]), .D(TxData[6]), .Z(n306) );
  AOI22CDNM1P U355 ( .A(TxData[0]), .B(TxData[1]), .C(TxData[1]), .D(TxData[0]), .Z(n298) );
  AOI22CDNM1P U356 ( .A(TxData[2]), .B(TxData[3]), .C(TxData[3]), .D(TxData[2]), .Z(n297) );
  N1M1P U357 ( .A(TxData[4]), .Z(n295) );
  AOI22CDNM1P U358 ( .A(TxData[5]), .B(n295), .C(n295), .D(TxData[5]), .Z(n296) );
  EN3M1P U359 ( .A(n298), .B(n297), .C(n296), .Z(n305) );
  AOI22CDNM1P U360 ( .A(TxData[15]), .B(TxData[16]), .C(TxData[16]), .D(
        TxData[15]), .Z(n302) );
  AOI22CDNM1P U361 ( .A(TxData[17]), .B(TxData[18]), .C(TxData[18]), .D(
        TxData[17]), .Z(n301) );
  N1M1P U362 ( .A(TxData[19]), .Z(n299) );
  AOI22CDNM1P U363 ( .A(TxData[23]), .B(n299), .C(n299), .D(TxData[23]), .Z(
        n300) );
  EN3M1P U364 ( .A(n302), .B(n301), .C(n300), .Z(n303) );
  EN3M1P U365 ( .A(TxData[22]), .B(TxData[14]), .C(n303), .Z(n304) );
  EN3M1P U366 ( .A(n306), .B(n305), .C(n304), .Z(n307) );
  EN3M1P U367 ( .A(n309), .B(n308), .C(n307), .Z(n316) );
  AOI22CDNM1P U368 ( .A(TxData[12]), .B(TxData[13]), .C(TxData[13]), .D(
        TxData[12]), .Z(n312) );
  AOI22CDNM1P U369 ( .A(TxData[8]), .B(TxData[9]), .C(TxData[9]), .D(TxData[8]), .Z(n311) );
  AOI22CDNM1P U370 ( .A(TxData[10]), .B(TxData[11]), .C(TxData[11]), .D(
        TxData[10]), .Z(n310) );
  EN3M1P U371 ( .A(n312), .B(n311), .C(n310), .Z(n313) );
  EN3M1P U372 ( .A(TxData[20]), .B(TxData[21]), .C(n313), .Z(n315) );
  ND2M1P U373 ( .A(n316), .B(n315), .Z(n314) );
  OAI211M1P U374 ( .A(n316), .B(n315), .C(n314), .D(n16), .Z(n317) );
  OAI21M1P U375 ( .A(n16), .B(n318), .C(n317), .Z(n157) );
  NR3M1P U376 ( .A(n273), .B(n329), .C(n327), .Z(n323) );
  NR2M1P U377 ( .A(n324), .B(n325), .Z(n322) );
  ND3M1P U378 ( .A(bitCount[3]), .B(n333), .C(n323), .Z(n321) );
  OAI22M1P U379 ( .A(n322), .B(n319), .C(n320), .D(n321), .Z(n28) );
  AOI22M1P U380 ( .A(bitCount[4]), .B(n322), .C(n321), .D(n320), .Z(n27) );
  AOI22M1P U381 ( .A(bitCount[3]), .B(n325), .C(n324), .D(n323), .Z(n326) );
  N1M1P U382 ( .A(n326), .Z(n26) );
  N1M1P U383 ( .A(n15), .Z(n339) );
  AOI21M1P U384 ( .A(n273), .B(n333), .C(n339), .Z(n330) );
  ND2M1P U385 ( .A(n333), .B(n329), .Z(n328) );
  AOI22M1P U386 ( .A(bitCount[0]), .B(n15), .C(n331), .D(n273), .Z(n23) );
  N1M1P U387 ( .A(n2), .Z(n343) );
  ND2M1P U388 ( .A(n344), .B(n343), .Z(n14) );
  NR2M1P U389 ( .A(n339), .B(n5), .Z(n332) );
  AOI211M1P U390 ( .A(n338), .B(n339), .C(n333), .D(n332), .Z(n12) );
  NR2M1P U391 ( .A(n7), .B(n93), .Z(n337) );
  N1M1P U392 ( .A(n11), .Z(n334) );
  OR3M1P U393 ( .A(n11), .B(n7), .C(n93), .Z(n336) );
  OAI211M1P U394 ( .A(n337), .B(n334), .C(n335), .D(n336), .Z(n10) );
  AO21CNM1P U395 ( .A(n9), .B(n336), .C(n335), .Z(n8) );
  AO211M1P U396 ( .A(n7), .B(n93), .C(Tx_Ready), .D(n337), .Z(n6) );
  ND3M1P U397 ( .A(n5), .B(n339), .C(n338), .Z(n342) );
endmodule

