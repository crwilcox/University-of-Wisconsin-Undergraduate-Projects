library verilog;
use verilog.vl_types.all;
entity prime_detector_behavioral_noglitch_tb is
    generic(
        SAMPLING_DELAY  : integer := 2
    );
end prime_detector_behavioral_noglitch_tb;
