library verilog;
use verilog.vl_types.all;
entity p8_exam1_solution is
end p8_exam1_solution;
